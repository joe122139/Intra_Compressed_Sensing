# Confidential Information of ARM, Inc.
# Use subject to ARM license.
# Copyright (c) 2017 ARM, Inc.

# ACI Version r1p1

# Reifier 4.0.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;

#name: High Density Two Port Register File RVT RVT Compiler | LOGIC0040LL 40nm Process 0.589um^2 Bit Cell
#version: r1p1
#comment: This is a memory instance
#configuration:  -activity_factor 50 -back_biasing off -bits 8 -bmux off -bus_notation on -check_instname on -diodes on -drive 6 -ema on -frequency 1.0 -instname rf_2p_hde -left_bus_delim "[" -mux 4 -mvt "" -name_case upper -power_type otc -prefix "" -pwr_gnd_rename vddpe:VDDPE,vddce:VDDCE,vsse:VSSE -retention on -right_bus_delim "]" -ser none -site_def off -top_layer m5-m10 -words 1024 -write_mask off -corners ff_1p21v_1p21v_125c,ff_1p21v_1p21v_m40c,ss_0p99v_0p99v_125c,ss_0p99v_0p99v_m40c,tt_1p10v_1p10v_25c
MACRO rf_2p_hde
  FOREIGN rf_2p_hde 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 110.215 BY 111.115 ;
  CLASS BLOCK ;
  PIN COLLDISN
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 53.21 0.0 53.35 0.25 ;
      LAYER M2 ;
      RECT 53.21 0.0 53.35 0.25 ;
      LAYER M3 ;
      RECT 53.21 0.0 53.35 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END COLLDISN
  PIN AA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 51.865 0.0 52.005 0.25 ;
      LAYER M2 ;
      RECT 51.865 0.0 52.005 0.25 ;
      LAYER M1 ;
      RECT 51.865 0.0 52.005 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[9]
  PIN AB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 58.25 0.0 58.39 0.25 ;
      LAYER M2 ;
      RECT 58.25 0.0 58.39 0.25 ;
      LAYER M3 ;
      RECT 58.25 0.0 58.39 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[9]
  PIN AA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 49.0 0.0 49.14 0.25 ;
      LAYER M2 ;
      RECT 49.0 0.0 49.14 0.25 ;
      LAYER M1 ;
      RECT 49.0 0.0 49.14 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[8]
  PIN AB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 61.075 0.0 61.215 0.25 ;
      LAYER M2 ;
      RECT 61.075 0.0 61.215 0.25 ;
      LAYER M3 ;
      RECT 61.075 0.0 61.215 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[8]
  PIN AA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 48.59 0.0 48.73 0.25 ;
      LAYER M2 ;
      RECT 48.59 0.0 48.73 0.25 ;
      LAYER M1 ;
      RECT 48.59 0.0 48.73 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[7]
  PIN AB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 61.485 0.0 61.625 0.25 ;
      LAYER M2 ;
      RECT 61.485 0.0 61.625 0.25 ;
      LAYER M3 ;
      RECT 61.485 0.0 61.625 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[7]
  PIN AA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 46.045 0.0 46.185 0.25 ;
      LAYER M2 ;
      RECT 46.045 0.0 46.185 0.25 ;
      LAYER M1 ;
      RECT 46.045 0.0 46.185 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[6]
  PIN AB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 64.045 0.0 64.185 0.25 ;
      LAYER M2 ;
      RECT 64.045 0.0 64.185 0.25 ;
      LAYER M3 ;
      RECT 64.045 0.0 64.185 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[6]
  PIN EMAA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.765 0.0 45.905 0.25 ;
      LAYER M2 ;
      RECT 45.765 0.0 45.905 0.25 ;
      LAYER M1 ;
      RECT 45.765 0.0 45.905 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAA[2]
  PIN EMAB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 64.325 0.0 64.465 0.25 ;
      LAYER M2 ;
      RECT 64.325 0.0 64.465 0.25 ;
      LAYER M3 ;
      RECT 64.325 0.0 64.465 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAB[2]
  PIN EMAA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 45.315 0.0 45.455 0.25 ;
      LAYER M3 ;
      RECT 45.315 0.0 45.455 0.25 ;
      LAYER M2 ;
      RECT 45.315 0.0 45.455 0.25 ;
      LAYER M1 ;
      RECT 45.315 0.0 45.455 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAA[1]
  PIN EMAB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 64.72 0.0 64.86 0.25 ;
      LAYER M2 ;
      RECT 64.72 0.0 64.86 0.25 ;
      LAYER M3 ;
      RECT 64.72 0.0 64.86 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAB[1]
  PIN AA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 45.03 0.0 45.17 0.25 ;
      LAYER M2 ;
      RECT 45.03 0.0 45.17 0.25 ;
      LAYER M1 ;
      RECT 45.03 0.0 45.17 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[5]
  PIN AB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 65.04 0.0 65.18 0.25 ;
      LAYER M2 ;
      RECT 65.04 0.0 65.18 0.25 ;
      LAYER M3 ;
      RECT 65.04 0.0 65.18 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[5]
  PIN EMAA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 44.545 0.0 44.685 0.25 ;
      LAYER M2 ;
      RECT 44.545 0.0 44.685 0.25 ;
      LAYER M1 ;
      RECT 44.545 0.0 44.685 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAA[0]
  PIN EMAB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 65.525 0.0 65.665 0.25 ;
      LAYER M2 ;
      RECT 65.525 0.0 65.665 0.25 ;
      LAYER M3 ;
      RECT 65.525 0.0 65.665 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END EMAB[0]
  PIN CENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 43.13 0.0 43.27 0.25 ;
      LAYER M2 ;
      RECT 43.13 0.0 43.27 0.25 ;
      LAYER M1 ;
      RECT 43.13 0.0 43.27 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CENA
  PIN CENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 66.95 0.0 67.09 0.25 ;
      LAYER M2 ;
      RECT 66.95 0.0 67.09 0.25 ;
      LAYER M3 ;
      RECT 66.95 0.0 67.09 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CENB
  PIN AA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 42.445 0.0 42.585 0.25 ;
      LAYER M2 ;
      RECT 42.445 0.0 42.585 0.25 ;
      LAYER M1 ;
      RECT 42.445 0.0 42.585 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[4]
  PIN AB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 67.63 0.0 67.77 0.25 ;
      LAYER M2 ;
      RECT 67.63 0.0 67.77 0.25 ;
      LAYER M3 ;
      RECT 67.63 0.0 67.77 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[4]
  PIN AA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 42.035 0.0 42.175 0.25 ;
      LAYER M2 ;
      RECT 42.035 0.0 42.175 0.25 ;
      LAYER M1 ;
      RECT 42.035 0.0 42.175 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[3]
  PIN AB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 68.04 0.0 68.18 0.25 ;
      LAYER M2 ;
      RECT 68.04 0.0 68.18 0.25 ;
      LAYER M3 ;
      RECT 68.04 0.0 68.18 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[3]
  PIN CLKA
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 40.65 0.0 40.79 0.25 ;
      LAYER M2 ;
      RECT 40.65 0.0 40.79 0.25 ;
      LAYER M1 ;
      RECT 40.65 0.0 40.79 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CLKA
  PIN CLKB
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 68.98 0.0 69.12 0.25 ;
      LAYER M2 ;
      RECT 68.98 0.0 69.12 0.25 ;
      LAYER M3 ;
      RECT 68.98 0.0 69.12 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END CLKB
  PIN AA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 39.165 0.0 39.305 0.25 ;
      LAYER M2 ;
      RECT 39.165 0.0 39.305 0.25 ;
      LAYER M1 ;
      RECT 39.165 0.0 39.305 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[2]
  PIN AB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 70.91 0.0 71.05 0.25 ;
      LAYER M2 ;
      RECT 70.91 0.0 71.05 0.25 ;
      LAYER M3 ;
      RECT 70.91 0.0 71.05 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[2]
  PIN AA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 38.755 0.0 38.895 0.25 ;
      LAYER M2 ;
      RECT 38.755 0.0 38.895 0.25 ;
      LAYER M1 ;
      RECT 38.755 0.0 38.895 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[1]
  PIN AB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 71.32 0.0 71.46 0.25 ;
      LAYER M2 ;
      RECT 71.32 0.0 71.46 0.25 ;
      LAYER M3 ;
      RECT 71.32 0.0 71.46 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[1]
  PIN AA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 35.89 0.0 36.03 0.25 ;
      LAYER M3 ;
      RECT 35.89 0.0 36.03 0.25 ;
      LAYER M2 ;
      RECT 35.89 0.0 36.03 0.25 ;
      LAYER M1 ;
      RECT 35.89 0.0 36.03 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AA[0]
  PIN AB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 74.145 0.0 74.285 0.25 ;
      LAYER M2 ;
      RECT 74.145 0.0 74.285 0.25 ;
      LAYER M3 ;
      RECT 74.145 0.0 74.285 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END AB[0]
  PIN RET1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 28.485 0.0 28.625 0.25 ;
      LAYER M2 ;
      RECT 28.485 0.0 28.625 0.25 ;
      LAYER M1 ;
      RECT 28.485 0.0 28.625 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END RET1N
  PIN DB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 84.855 0.0 84.995 0.25 ;
      LAYER M2 ;
      RECT 84.855 0.0 84.995 0.25 ;
      LAYER M3 ;
      RECT 84.855 0.0 84.995 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[4]
  PIN DB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 25.22 0.0 25.36 0.25 ;
      LAYER M2 ;
      RECT 25.22 0.0 25.36 0.25 ;
      LAYER M1 ;
      RECT 25.22 0.0 25.36 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[3]
  PIN QA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 87.345 0.0 87.485 0.25 ;
      LAYER M2 ;
      RECT 87.345 0.0 87.485 0.25 ;
      LAYER M3 ;
      RECT 87.345 0.0 87.485 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[4]
  PIN QA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 22.73 0.0 22.87 0.25 ;
      LAYER M2 ;
      RECT 22.73 0.0 22.87 0.25 ;
      LAYER M1 ;
      RECT 22.73 0.0 22.87 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[3]
  PIN DB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 91.055 0.0 91.195 0.25 ;
      LAYER M2 ;
      RECT 91.055 0.0 91.195 0.25 ;
      LAYER M3 ;
      RECT 91.055 0.0 91.195 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[5]
  PIN DB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 19.02 0.0 19.16 0.25 ;
      LAYER M2 ;
      RECT 19.02 0.0 19.16 0.25 ;
      LAYER M1 ;
      RECT 19.02 0.0 19.16 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[2]
  PIN QA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 93.545 0.0 93.685 0.25 ;
      LAYER M2 ;
      RECT 93.545 0.0 93.685 0.25 ;
      LAYER M3 ;
      RECT 93.545 0.0 93.685 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[5]
  PIN QA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 16.53 0.0 16.67 0.25 ;
      LAYER M2 ;
      RECT 16.53 0.0 16.67 0.25 ;
      LAYER M1 ;
      RECT 16.53 0.0 16.67 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[2]
  PIN DB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 97.255 0.0 97.395 0.25 ;
      LAYER M2 ;
      RECT 97.255 0.0 97.395 0.25 ;
      LAYER M3 ;
      RECT 97.255 0.0 97.395 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[6]
  PIN DB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 12.82 0.0 12.96 0.25 ;
      LAYER M2 ;
      RECT 12.82 0.0 12.96 0.25 ;
      LAYER M1 ;
      RECT 12.82 0.0 12.96 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[1]
  PIN QA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 99.745 0.0 99.885 0.25 ;
      LAYER M2 ;
      RECT 99.745 0.0 99.885 0.25 ;
      LAYER M3 ;
      RECT 99.745 0.0 99.885 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[6]
  PIN QA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 10.33 0.0 10.47 0.25 ;
      LAYER M2 ;
      RECT 10.33 0.0 10.47 0.25 ;
      LAYER M1 ;
      RECT 10.33 0.0 10.47 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[1]
  PIN DB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 103.455 0.0 103.595 0.25 ;
      LAYER M2 ;
      RECT 103.455 0.0 103.595 0.25 ;
      LAYER M3 ;
      RECT 103.455 0.0 103.595 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[7]
  PIN DB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 6.62 0.0 6.76 0.25 ;
      LAYER M2 ;
      RECT 6.62 0.0 6.76 0.25 ;
      LAYER M1 ;
      RECT 6.62 0.0 6.76 0.25 ;
      END
    ANTENNAGATEAREA 0.0114 ;
    ANTENNADIFFAREA 0.035 ;
    END DB[0]
  PIN QA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT 105.945 0.0 106.085 0.25 ;
      LAYER M2 ;
      RECT 105.945 0.0 106.085 0.25 ;
      LAYER M3 ;
      RECT 105.945 0.0 106.085 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[7]
  PIN QA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M3 ;
      RECT 4.13 0.0 4.27 0.25 ;
      LAYER M2 ;
      RECT 4.13 0.0 4.27 0.25 ;
      LAYER M1 ;
      RECT 4.13 0.0 4.27 0.25 ;
      END
    ANTENNADIFFAREA 0.035 ;
    END QA[0]
  PIN VDDPE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.72 0.0 0.86 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 3.66 0.0 3.94 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 6.76 0.0 7.04 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 9.86 0.0 10.14 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 12.96 0.0 13.24 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 16.06 0.0 16.34 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 19.16 0.0 19.44 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 22.26 0.0 22.54 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.36 0.0 25.64 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 25.8 0.0 26.01 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 28.12 0.0 28.4 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 30.915 0.0 31.195 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 35.105 0.0 35.385 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 36.505 0.0 36.785 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 39.3 0.0 39.58 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 40.695 0.0 40.975 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 42.095 0.0 42.375 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 46.285 0.0 46.565 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 47.68 0.0 47.96 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 51.875 0.0 52.155 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 53.27 0.0 53.55 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 56.765 0.0 57.045 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 58.16 0.0 58.44 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 62.35 0.0 62.63 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 63.75 0.0 64.03 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 67.94 0.0 68.22 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 69.335 0.0 69.615 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 70.735 0.0 71.015 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 73.535 0.0 73.815 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 74.935 0.0 75.215 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 79.12 0.0 79.4 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 81.915 0.0 82.195 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 84.205 0.0 84.415 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 84.575 0.0 84.855 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 87.675 0.0 87.955 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 90.775 0.0 91.055 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 93.875 0.0 94.155 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 96.975 0.0 97.255 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.075 0.0 100.355 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 103.175 0.0 103.455 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 106.275 0.0 106.555 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 109.355 0.0 109.495 111.115 ;
      END
    END VDDPE
  PIN VDDCE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.16 0.0 0.3 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 1.66 0.0 1.94 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 4.76 0.0 5.04 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 7.86 0.0 8.14 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 10.96 0.0 11.24 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 14.06 0.0 14.34 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 17.16 0.0 17.44 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 20.26 0.0 20.54 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 23.36 0.0 23.64 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 26.5 0.0 26.71 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 32.31 0.0 32.59 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 33.71 0.0 33.99 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.9 0.0 38.18 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 43.49 0.0 43.77 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 44.89 0.0 45.17 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 49.08 0.0 49.36 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 50.475 0.0 50.755 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 54.67 0.0 54.95 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 55.365 0.0 55.645 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 59.56 0.0 59.84 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 60.955 0.0 61.235 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 65.145 0.0 65.425 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 66.545 0.0 66.825 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 72.135 0.0 72.415 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 76.325 0.0 76.605 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 77.72 0.0 78.0 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 83.505 0.0 83.715 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 86.575 0.0 86.855 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 89.675 0.0 89.955 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 92.775 0.0 93.055 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 95.875 0.0 96.155 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 98.975 0.0 99.255 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 102.075 0.0 102.355 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 105.175 0.0 105.455 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 108.275 0.0 108.555 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 109.915 0.0 110.055 111.115 ;
      END
    END VDDCE
  PIN VSSE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.44 0.0 0.58 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 3.005 0.0 3.285 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 6.105 0.0 6.385 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 9.205 0.0 9.485 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 12.305 0.0 12.585 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 15.405 0.0 15.685 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 18.505 0.0 18.785 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 21.605 0.0 21.885 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 24.705 0.0 24.985 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 26.15 0.0 26.36 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 27.42 0.0 27.7 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 28.82 0.0 29.1 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 31.615 0.0 31.895 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 33.01 0.0 33.29 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 34.41 0.0 34.69 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 37.205 0.0 37.485 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 38.6 0.0 38.88 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 39.995 0.0 40.275 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 42.79 0.0 43.07 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 44.19 0.0 44.47 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 45.585 0.0 45.865 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 48.38 0.0 48.66 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 49.78 0.0 50.06 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 53.97 0.0 54.25 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 56.065 0.0 56.345 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 60.26 0.0 60.54 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 61.655 0.0 61.935 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 64.445 0.0 64.725 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 65.845 0.0 66.125 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 67.24 0.0 67.52 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 70.035 0.0 70.315 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 71.435 0.0 71.715 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 72.835 0.0 73.115 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 75.635 0.0 75.915 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 77.02 0.0 77.3 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 78.42 0.0 78.7 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 81.215 0.0 81.495 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 82.615 0.0 82.895 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 83.855 0.0 84.065 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 85.23 0.0 85.51 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 88.33 0.0 88.61 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 91.43 0.0 91.71 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 94.53 0.0 94.81 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 97.63 0.0 97.91 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 100.73 0.0 101.01 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 103.83 0.0 104.11 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 106.93 0.0 107.21 111.115 ;
      END
    PORT
      LAYER M4 ;
      RECT 109.635 0.0 109.775 111.115 ;
      END
    END VSSE
  OBS
    #otc obstructions
    LAYER M1 DESIGNRULEWIDTH 0.07 ;
    RECT 106.225 0.0 110.215 0.32 ;
    RECT 103.735 0.0 105.805 0.32 ;
    RECT 100.025 0.0 103.315 0.32 ;
    RECT 97.535 0.0 99.605 0.32 ;
    RECT 93.825 0.0 97.115 0.32 ;
    RECT 91.335 0.0 93.405 0.32 ;
    RECT 87.625 0.0 90.915 0.32 ;
    RECT 85.135 0.0 87.205 0.32 ;
    RECT 74.425 0.0 84.715 0.32 ;
    RECT 71.6 0.0 74.005 0.32 ;
    RECT 69.26 0.0 70.77 0.32 ;
    RECT 68.32 0.0 68.84 0.32 ;
    RECT 67.23 0.0 67.49 0.32 ;
    RECT 65.805 0.0 66.81 0.32 ;
    RECT 61.765 0.0 63.905 0.32 ;
    RECT 58.53 0.0 60.935 0.32 ;
    RECT 53.49 0.0 58.11 0.32 ;
    RECT 52.145 0.0 53.07 0.32 ;
    RECT 49.28 0.0 51.725 0.32 ;
    RECT 46.325 0.0 48.45 0.32 ;
    RECT 43.41 0.0 44.405 0.32 ;
    RECT 42.725 0.0 42.99 0.32 ;
    RECT 40.93 0.0 41.895 0.32 ;
    RECT 39.445 0.0 40.51 0.32 ;
    RECT 36.17 0.0 38.615 0.32 ;
    RECT 28.765 0.0 35.75 0.32 ;
    RECT 25.5 0.0 28.345 0.32 ;
    RECT 23.01 0.0 25.08 0.32 ;
    RECT 19.3 0.0 22.59 0.32 ;
    RECT 16.81 0.0 18.88 0.32 ;
    RECT 13.1 0.0 16.39 0.32 ;
    RECT 10.61 0.0 12.68 0.32 ;
    RECT 6.9 0.0 10.19 0.32 ;
    RECT 4.41 0.0 6.48 0.32 ;
    RECT 0.0 0.0 3.99 0.32 ;
    RECT 0.0 0.32 110.215 111.115 ;
    LAYER V1 ;
    RECT 0.0 0.0 110.215 111.115 ;
    LAYER M2 DESIGNRULEWIDTH 0.07 ;
    RECT 106.225 0.0 110.215 0.32 ;
    RECT 103.735 0.0 105.805 0.32 ;
    RECT 100.025 0.0 103.315 0.32 ;
    RECT 97.535 0.0 99.605 0.32 ;
    RECT 93.825 0.0 97.115 0.32 ;
    RECT 91.335 0.0 93.405 0.32 ;
    RECT 87.625 0.0 90.915 0.32 ;
    RECT 85.135 0.0 87.205 0.32 ;
    RECT 74.425 0.0 84.715 0.32 ;
    RECT 71.6 0.0 74.005 0.32 ;
    RECT 69.26 0.0 70.77 0.32 ;
    RECT 68.32 0.0 68.84 0.32 ;
    RECT 67.23 0.0 67.49 0.32 ;
    RECT 65.805 0.0 66.81 0.32 ;
    RECT 61.765 0.0 63.905 0.32 ;
    RECT 58.53 0.0 60.935 0.32 ;
    RECT 53.49 0.0 58.11 0.32 ;
    RECT 52.145 0.0 53.07 0.32 ;
    RECT 49.28 0.0 51.725 0.32 ;
    RECT 46.325 0.0 48.45 0.32 ;
    RECT 43.41 0.0 44.405 0.32 ;
    RECT 42.725 0.0 42.99 0.32 ;
    RECT 40.93 0.0 41.895 0.32 ;
    RECT 39.445 0.0 40.51 0.32 ;
    RECT 36.17 0.0 38.615 0.32 ;
    RECT 28.765 0.0 35.75 0.32 ;
    RECT 25.5 0.0 28.345 0.32 ;
    RECT 23.01 0.0 25.08 0.32 ;
    RECT 19.3 0.0 22.59 0.32 ;
    RECT 16.81 0.0 18.88 0.32 ;
    RECT 13.1 0.0 16.39 0.32 ;
    RECT 10.61 0.0 12.68 0.32 ;
    RECT 6.9 0.0 10.19 0.32 ;
    RECT 4.41 0.0 6.48 0.32 ;
    RECT 0.0 0.0 3.99 0.32 ;
    RECT 0.0 0.32 110.215 111.115 ;
    LAYER V2 ;
    RECT 0.0 0.0 110.215 111.115 ;
    LAYER M3 DESIGNRULEWIDTH 0.07 ;
    RECT 106.225 0.0 110.215 0.32 ;
    RECT 103.735 0.0 105.805 0.32 ;
    RECT 100.025 0.0 103.315 0.32 ;
    RECT 97.535 0.0 99.605 0.32 ;
    RECT 93.825 0.0 97.115 0.32 ;
    RECT 91.335 0.0 93.405 0.32 ;
    RECT 87.625 0.0 90.915 0.32 ;
    RECT 85.135 0.0 87.205 0.32 ;
    RECT 74.425 0.0 84.715 0.32 ;
    RECT 71.6 0.0 74.005 0.32 ;
    RECT 69.26 0.0 70.77 0.32 ;
    RECT 68.32 0.0 68.84 0.32 ;
    RECT 67.23 0.0 67.49 0.32 ;
    RECT 65.805 0.0 66.81 0.32 ;
    RECT 61.765 0.0 63.905 0.32 ;
    RECT 58.53 0.0 60.935 0.32 ;
    RECT 53.49 0.0 58.11 0.32 ;
    RECT 52.145 0.0 53.07 0.32 ;
    RECT 49.28 0.0 51.725 0.32 ;
    RECT 46.325 0.0 48.45 0.32 ;
    RECT 43.41 0.0 44.405 0.32 ;
    RECT 42.725 0.0 42.99 0.32 ;
    RECT 40.93 0.0 41.895 0.32 ;
    RECT 39.445 0.0 40.51 0.32 ;
    RECT 36.17 0.0 38.615 0.32 ;
    RECT 28.765 0.0 35.75 0.32 ;
    RECT 25.5 0.0 28.345 0.32 ;
    RECT 23.01 0.0 25.08 0.32 ;
    RECT 19.3 0.0 22.59 0.32 ;
    RECT 16.81 0.0 18.88 0.32 ;
    RECT 13.1 0.0 16.39 0.32 ;
    RECT 10.61 0.0 12.68 0.32 ;
    RECT 6.9 0.0 10.19 0.32 ;
    RECT 4.41 0.0 6.48 0.32 ;
    RECT 0.0 0.0 3.99 0.32 ;
    RECT 0.0 0.32 110.215 111.115 ;
    LAYER V3 ;
    RECT 0.0 0.0 110.215 111.115 ;
    LAYER V3 ;
    RECT 75.67 0.645 75.88 0.715 ;
    RECT 34.445 0.645 34.655 0.715 ;
    RECT 26.15 0.645 26.36 0.715 ;
    RECT 79.855 0.645 80.065 0.715 ;
    RECT 74.27 0.645 74.48 0.715 ;
    RECT 47.715 9.475 47.925 9.685 ;
    RECT 47.715 8.09 47.925 8.16 ;
    RECT 47.715 3.26 47.925 3.33 ;
    RECT 72.87 7.09 73.08 7.16 ;
    RECT 72.87 3.65 73.08 3.72 ;
    RECT 72.87 1.375 73.08 1.585 ;
    RECT 47.715 0.885 47.925 1.095 ;
    RECT 30.25 2.86 30.46 2.93 ;
    RECT 68.675 0.645 68.885 0.715 ;
    RECT 63.085 0.645 63.295 0.715 ;
    RECT 57.5 0.645 57.71 0.715 ;
    RECT 46.32 4.72 46.53 4.79 ;
    RECT 71.47 7.09 71.68 7.16 ;
    RECT 46.32 2.01 46.53 2.08 ;
    RECT 71.47 3.65 71.68 3.72 ;
    RECT 71.47 1.375 71.68 1.585 ;
    RECT 42.13 4.72 42.34 4.79 ;
    RECT 70.07 7.09 70.28 7.16 ;
    RECT 28.855 7.09 29.065 7.16 ;
    RECT 52.61 0.645 52.82 0.715 ;
    RECT 47.02 0.645 47.23 0.715 ;
    RECT 41.43 0.645 41.64 0.715 ;
    RECT 35.84 0.645 36.05 0.715 ;
    RECT 42.13 2.01 42.34 2.08 ;
    RECT 70.07 3.65 70.28 3.72 ;
    RECT 70.07 1.375 70.28 1.585 ;
    RECT 40.73 4.72 40.94 4.79 ;
    RECT 40.73 2.01 40.94 2.08 ;
    RECT 39.335 4.72 39.545 4.79 ;
    RECT 28.855 3.65 29.065 3.72 ;
    RECT 39.335 2.01 39.545 2.08 ;
    RECT 28.855 1.375 29.065 1.585 ;
    RECT 27.455 7.09 27.665 7.16 ;
    RECT 68.675 2.86 68.885 2.93 ;
    RECT 27.455 3.65 27.665 3.72 ;
    RECT 27.455 1.375 27.665 1.585 ;
    RECT 30.25 0.645 30.46 0.715 ;
    RECT 36.54 4.72 36.75 4.79 ;
    RECT 36.54 2.01 36.75 2.08 ;
    RECT 35.14 4.72 35.35 4.79 ;
    RECT 35.14 2.01 35.35 2.08 ;
    RECT 67.275 7.09 67.485 7.16 ;
    RECT 67.275 3.65 67.485 3.72 ;
    RECT 67.275 1.375 67.485 1.585 ;
    RECT 65.88 7.09 66.09 7.16 ;
    RECT 65.88 3.65 66.09 3.72 ;
    RECT 65.88 1.375 66.09 1.585 ;
    RECT 64.48 7.09 64.69 7.16 ;
    RECT 64.48 3.65 64.69 3.72 ;
    RECT 30.95 4.72 31.16 4.79 ;
    RECT 30.95 2.01 31.16 2.08 ;
    RECT 64.48 1.375 64.69 1.585 ;
    RECT 63.085 2.86 63.295 2.93 ;
    RECT 28.155 4.72 28.365 4.79 ;
    RECT 28.155 2.01 28.365 2.08 ;
    RECT 25.8 9.475 26.01 9.685 ;
    RECT 61.69 7.09 61.9 7.16 ;
    RECT 61.69 3.65 61.9 3.72 ;
    RECT 61.69 1.375 61.9 1.585 ;
    RECT 25.8 8.09 26.01 8.16 ;
    RECT 25.8 3.26 26.01 3.33 ;
    RECT 25.8 0.885 26.01 1.095 ;
    RECT 60.295 7.09 60.505 7.16 ;
    RECT 60.295 3.65 60.505 3.72 ;
    RECT 60.295 1.375 60.505 1.585 ;
    RECT 57.5 2.86 57.71 2.93 ;
    RECT 80.55 9.3 80.76 9.37 ;
    RECT 77.755 9.1 77.965 9.17 ;
    RECT 76.36 9.1 76.57 9.17 ;
    RECT 72.17 9.1 72.38 9.17 ;
    RECT 66.58 9.1 66.79 9.17 ;
    RECT 65.18 9.1 65.39 9.17 ;
    RECT 60.99 9.1 61.2 9.17 ;
    RECT 56.1 7.09 56.31 7.16 ;
    RECT 56.1 3.65 56.31 3.72 ;
    RECT 56.1 1.375 56.31 1.585 ;
    RECT 55.4 9.1 55.61 9.17 ;
    RECT 54.705 9.1 54.915 9.17 ;
    RECT 49.115 9.1 49.325 9.17 ;
    RECT 44.925 9.1 45.135 9.17 ;
    RECT 43.525 9.1 43.735 9.17 ;
    RECT 37.935 9.1 38.145 9.17 ;
    RECT 33.745 9.1 33.955 9.17 ;
    RECT 32.345 9.1 32.555 9.17 ;
    RECT 34.415 0.245 34.675 0.315 ;
    RECT 35.925 0.06 35.995 0.27 ;
    RECT 45.35 0.06 45.42 0.27 ;
    RECT 74.665 0.06 74.735 0.27 ;
    RECT 75.635 0.245 75.895 0.315 ;
    RECT 84.205 9.475 84.415 9.685 ;
    RECT 82.65 6.31 82.86 6.38 ;
    RECT 81.25 6.31 81.46 6.38 ;
    RECT 54.005 7.09 54.215 7.16 ;
    RECT 54.005 3.65 54.215 3.72 ;
    RECT 54.005 1.375 54.215 1.585 ;
    RECT 29.555 9.3 29.765 9.37 ;
    RECT 84.205 8.09 84.415 8.16 ;
    RECT 84.205 3.26 84.415 3.33 ;
    RECT 78.455 6.31 78.665 6.38 ;
    RECT 84.205 0.885 84.415 1.095 ;
    RECT 81.95 4.72 82.16 4.79 ;
    RECT 77.055 6.31 77.265 6.38 ;
    RECT 81.95 2.01 82.16 2.08 ;
    RECT 75.67 2.86 75.88 2.93 ;
    RECT 52.61 2.86 52.82 2.93 ;
    RECT 72.87 6.31 73.08 6.38 ;
    RECT 71.47 6.31 71.68 6.38 ;
    RECT 70.07 6.31 70.28 6.38 ;
    RECT 49.815 7.09 50.025 7.16 ;
    RECT 49.815 3.65 50.025 3.72 ;
    RECT 49.815 1.375 50.025 1.585 ;
    RECT 79.155 4.72 79.365 4.79 ;
    RECT 79.155 2.01 79.365 2.08 ;
    RECT 67.275 6.31 67.485 6.38 ;
    RECT 65.88 6.31 66.09 6.38 ;
    RECT 64.48 6.31 64.69 6.38 ;
    RECT 48.415 7.09 48.625 7.16 ;
    RECT 48.415 3.65 48.625 3.72 ;
    RECT 61.69 6.31 61.9 6.38 ;
    RECT 48.415 1.375 48.625 1.585 ;
    RECT 47.02 2.86 47.23 2.93 ;
    RECT 60.295 6.31 60.505 6.38 ;
    RECT 45.62 7.09 45.83 7.16 ;
    RECT 56.1 6.31 56.31 6.38 ;
    RECT 45.62 3.65 45.83 3.86 ;
    RECT 54.005 6.31 54.215 6.38 ;
    RECT 45.62 1.375 45.83 1.585 ;
    RECT 74.97 4.72 75.18 4.79 ;
    RECT 44.225 7.09 44.435 7.16 ;
    RECT 74.97 2.01 75.18 2.08 ;
    RECT 44.225 3.65 44.435 3.72 ;
    RECT 73.57 4.72 73.78 4.79 ;
    RECT 73.57 2.01 73.78 2.08 ;
    RECT 27.43 9.83 27.69 9.9 ;
    RECT 28.83 9.83 29.09 9.9 ;
    RECT 31.625 9.83 31.885 9.9 ;
    RECT 33.025 9.83 33.285 9.9 ;
    RECT 37.22 9.83 37.475 9.9 ;
    RECT 38.615 9.83 38.875 9.9 ;
    RECT 40.01 9.83 40.27 9.9 ;
    RECT 41.395 7.105 41.67 7.175 ;
    RECT 42.805 9.83 43.065 9.9 ;
    RECT 44.205 9.83 44.465 9.9 ;
    RECT 45.6 9.83 45.86 9.9 ;
    RECT 48.385 9.83 48.655 9.9 ;
    RECT 49.78 9.83 50.05 9.9 ;
    RECT 52.575 7.105 52.845 7.175 ;
    RECT 53.725 2.01 53.795 2.08 ;
    RECT 53.725 4.725 53.795 4.795 ;
    RECT 53.97 9.83 54.245 9.9 ;
    RECT 56.07 9.83 56.34 9.9 ;
    RECT 60.26 9.83 60.525 9.9 ;
    RECT 61.655 9.83 61.92 9.9 ;
    RECT 64.46 9.83 64.725 9.9 ;
    RECT 65.86 9.83 66.12 9.9 ;
    RECT 67.245 9.83 67.505 9.9 ;
    RECT 68.645 7.105 68.915 7.175 ;
    RECT 70.04 9.83 70.3 9.9 ;
    RECT 71.44 9.83 71.705 9.9 ;
    RECT 72.85 9.83 73.105 9.9 ;
    RECT 77.025 9.83 77.285 9.9 ;
    RECT 77.725 9.3 78.0 9.37 ;
    RECT 78.425 9.83 78.685 9.9 ;
    RECT 81.22 9.83 81.49 9.9 ;
    RECT 82.615 9.83 82.89 9.9 ;
    RECT 49.815 6.31 50.025 6.38 ;
    RECT 48.415 6.31 48.625 6.38 ;
    RECT 44.225 1.375 44.435 1.585 ;
    RECT 45.62 6.31 45.83 6.38 ;
    RECT 44.225 6.31 44.435 6.38 ;
    RECT 42.825 7.09 43.035 7.16 ;
    RECT 42.825 3.65 43.035 3.72 ;
    RECT 42.825 6.31 43.035 6.38 ;
    RECT 70.77 4.72 70.98 4.79 ;
    RECT 42.825 1.375 43.035 1.585 ;
    RECT 70.77 2.01 70.98 2.08 ;
    RECT 69.37 4.72 69.58 4.79 ;
    RECT 69.37 2.01 69.58 2.08 ;
    RECT 67.975 4.72 68.185 4.79 ;
    RECT 67.975 2.01 68.185 2.08 ;
    RECT 40.03 6.31 40.24 6.38 ;
    RECT 38.635 6.31 38.845 6.38 ;
    RECT 37.24 6.31 37.45 6.38 ;
    RECT 37.24 4.875 37.45 4.945 ;
    RECT 63.785 4.72 63.995 4.79 ;
    RECT 63.785 2.01 63.995 2.08 ;
    RECT 82.65 7.09 82.86 7.16 ;
    RECT 82.65 3.65 82.86 3.72 ;
    RECT 82.65 1.375 82.86 1.585 ;
    RECT 41.43 2.86 41.64 2.93 ;
    RECT 62.385 9.475 62.595 9.685 ;
    RECT 62.385 8.09 62.595 8.16 ;
    RECT 40.03 7.09 40.24 7.16 ;
    RECT 40.03 3.65 40.24 3.72 ;
    RECT 40.03 1.375 40.24 1.585 ;
    RECT 38.635 7.09 38.845 7.16 ;
    RECT 38.635 3.65 38.845 3.72 ;
    RECT 34.445 2.86 34.655 2.93 ;
    RECT 33.045 6.31 33.255 6.38 ;
    RECT 31.65 6.31 31.86 6.38 ;
    RECT 28.855 6.31 29.065 6.38 ;
    RECT 62.385 3.26 62.595 3.33 ;
    RECT 62.385 2.17 62.595 2.24 ;
    RECT 81.25 7.09 81.46 7.16 ;
    RECT 81.25 3.65 81.46 3.72 ;
    RECT 81.25 1.375 81.46 1.585 ;
    RECT 79.855 2.86 80.065 2.93 ;
    RECT 62.385 0.885 62.595 1.095 ;
    RECT 38.635 1.375 38.845 1.585 ;
    RECT 78.455 7.09 78.665 7.16 ;
    RECT 78.455 3.65 78.665 3.72 ;
    RECT 37.24 7.09 37.45 7.16 ;
    RECT 78.455 1.375 78.665 1.585 ;
    RECT 37.24 3.65 37.45 3.72 ;
    RECT 37.24 1.375 37.45 1.585 ;
    RECT 27.455 6.31 27.665 6.38 ;
    RECT 58.195 4.72 58.405 4.79 ;
    RECT 58.195 2.01 58.405 2.08 ;
    RECT 56.8 4.72 57.01 4.79 ;
    RECT 56.8 2.01 57.01 2.08 ;
    RECT 35.84 2.86 36.05 2.93 ;
    RECT 33.045 7.09 33.255 7.16 ;
    RECT 33.045 3.65 33.255 3.72 ;
    RECT 33.045 1.375 33.255 1.585 ;
    RECT 83.855 0.645 84.065 0.715 ;
    RECT 78.455 0.245 78.665 0.315 ;
    RECT 77.055 7.09 77.265 7.16 ;
    RECT 53.71 8.1 53.78 8.17 ;
    RECT 77.055 3.65 77.265 3.72 ;
    RECT 53.71 3.27 53.78 3.34 ;
    RECT 77.055 1.375 77.265 1.585 ;
    RECT 53.305 4.72 53.515 4.79 ;
    RECT 53.305 2.01 53.515 2.08 ;
    RECT 51.91 4.72 52.12 4.79 ;
    RECT 31.65 7.09 31.86 7.16 ;
    RECT 51.91 2.01 52.12 2.08 ;
    RECT 74.27 2.86 74.48 2.93 ;
    RECT 31.65 3.65 31.86 3.72 ;
    RECT 31.65 1.375 31.86 1.585 ;
    RECT 96.57 110.86 96.78 110.93 ;
    RECT 93.47 110.86 93.68 110.93 ;
    RECT 90.37 110.86 90.58 110.93 ;
    RECT 102.77 110.86 102.98 110.93 ;
    RECT 99.67 110.86 99.88 110.93 ;
    RECT 108.97 110.86 109.18 110.93 ;
    RECT 105.87 110.86 106.08 110.93 ;
    RECT 87.27 110.86 87.48 110.93 ;
    RECT 89.71 60.132 89.92 60.202 ;
    RECT 88.365 60.385 88.575 60.455 ;
    RECT 89.71 109.758 89.92 109.828 ;
    RECT 89.71 10.752 89.92 10.822 ;
    RECT 88.365 109.505 88.575 109.575 ;
    RECT 88.365 11.005 88.575 11.075 ;
    RECT 89.71 110.315 89.92 110.525 ;
    RECT 89.71 10.055 89.92 10.265 ;
    RECT 102.11 60.132 102.32 60.202 ;
    RECT 100.765 60.385 100.975 60.455 ;
    RECT 102.11 109.758 102.32 109.828 ;
    RECT 102.11 10.752 102.32 10.822 ;
    RECT 100.765 109.505 100.975 109.575 ;
    RECT 100.765 11.005 100.975 11.075 ;
    RECT 102.11 110.315 102.32 110.525 ;
    RECT 102.11 10.055 102.32 10.265 ;
    RECT 99.01 60.132 99.22 60.202 ;
    RECT 97.665 60.385 97.875 60.455 ;
    RECT 99.01 109.758 99.22 109.828 ;
    RECT 99.01 10.752 99.22 10.822 ;
    RECT 97.665 109.505 97.875 109.575 ;
    RECT 97.665 11.005 97.875 11.075 ;
    RECT 99.01 110.315 99.22 110.525 ;
    RECT 99.01 10.055 99.22 10.265 ;
    RECT 95.91 60.132 96.12 60.202 ;
    RECT 94.565 60.385 94.775 60.455 ;
    RECT 95.91 109.758 96.12 109.828 ;
    RECT 95.91 10.752 96.12 10.822 ;
    RECT 94.565 109.505 94.775 109.575 ;
    RECT 94.565 11.005 94.775 11.075 ;
    RECT 95.91 110.315 96.12 110.525 ;
    RECT 95.91 10.055 96.12 10.265 ;
    RECT 92.81 60.132 93.02 60.202 ;
    RECT 91.465 60.385 91.675 60.455 ;
    RECT 92.81 109.758 93.02 109.828 ;
    RECT 92.81 10.752 93.02 10.822 ;
    RECT 91.465 109.505 91.675 109.575 ;
    RECT 91.465 11.005 91.675 11.075 ;
    RECT 92.81 110.315 93.02 110.525 ;
    RECT 92.81 10.055 93.02 10.265 ;
    RECT 105.21 60.132 105.42 60.202 ;
    RECT 103.865 60.385 104.075 60.455 ;
    RECT 105.21 109.758 105.42 109.828 ;
    RECT 105.21 10.752 105.42 10.822 ;
    RECT 103.865 109.505 104.075 109.575 ;
    RECT 103.865 11.005 104.075 11.075 ;
    RECT 105.21 110.315 105.42 110.525 ;
    RECT 105.21 10.055 105.42 10.265 ;
    RECT 86.61 60.132 86.82 60.202 ;
    RECT 85.265 60.385 85.475 60.455 ;
    RECT 86.61 109.758 86.82 109.828 ;
    RECT 86.61 10.752 86.82 10.822 ;
    RECT 85.265 109.505 85.475 109.575 ;
    RECT 85.265 11.005 85.475 11.075 ;
    RECT 86.61 110.315 86.82 110.525 ;
    RECT 86.61 10.055 86.82 10.265 ;
    RECT 108.31 60.132 108.52 60.202 ;
    RECT 106.965 60.385 107.175 60.455 ;
    RECT 108.31 109.758 108.52 109.828 ;
    RECT 108.31 10.752 108.52 10.822 ;
    RECT 106.965 109.505 107.175 109.575 ;
    RECT 106.965 11.005 107.175 11.075 ;
    RECT 108.31 110.315 108.52 110.525 ;
    RECT 108.31 10.055 108.52 10.265 ;
    RECT 83.855 110.815 84.065 111.025 ;
    RECT 75.67 110.815 75.88 111.025 ;
    RECT 34.445 110.815 34.655 111.025 ;
    RECT 26.15 110.815 26.36 111.025 ;
    RECT 52.61 110.815 52.82 111.025 ;
    RECT 47.02 110.815 47.23 111.025 ;
    RECT 79.855 110.815 80.065 111.025 ;
    RECT 41.43 110.815 41.64 111.025 ;
    RECT 74.27 110.815 74.48 111.025 ;
    RECT 35.84 110.815 36.05 111.025 ;
    RECT 30.25 110.815 30.46 111.025 ;
    RECT 68.675 110.815 68.885 111.025 ;
    RECT 78.455 11.005 78.665 11.075 ;
    RECT 77.055 11.005 77.265 11.075 ;
    RECT 72.87 11.005 73.08 11.075 ;
    RECT 71.47 11.005 71.68 11.075 ;
    RECT 70.07 11.005 70.28 11.075 ;
    RECT 67.275 11.005 67.485 11.075 ;
    RECT 65.88 11.005 66.09 11.075 ;
    RECT 64.48 11.005 64.69 11.075 ;
    RECT 61.69 11.005 61.9 11.075 ;
    RECT 60.295 11.005 60.505 11.075 ;
    RECT 56.1 11.005 56.31 11.075 ;
    RECT 54.005 11.005 54.215 11.075 ;
    RECT 49.815 11.005 50.025 11.075 ;
    RECT 29.525 11.625 30.74 11.695 ;
    RECT 29.525 12.385 30.74 12.455 ;
    RECT 29.525 13.145 30.74 13.215 ;
    RECT 29.525 13.905 30.74 13.975 ;
    RECT 29.525 14.665 30.74 14.735 ;
    RECT 29.525 15.425 30.74 15.495 ;
    RECT 29.525 16.185 30.74 16.255 ;
    RECT 29.525 16.945 30.74 17.015 ;
    RECT 29.525 17.705 30.74 17.775 ;
    RECT 29.525 18.465 30.74 18.535 ;
    RECT 29.525 19.225 30.74 19.295 ;
    RECT 29.525 19.985 30.74 20.055 ;
    RECT 29.525 20.745 30.74 20.815 ;
    RECT 29.525 21.505 30.74 21.575 ;
    RECT 29.525 22.265 30.74 22.335 ;
    RECT 29.525 23.025 30.74 23.095 ;
    RECT 53.975 11.625 54.245 11.695 ;
    RECT 53.975 12.385 54.245 12.455 ;
    RECT 53.975 13.145 54.245 13.215 ;
    RECT 53.975 13.905 54.245 13.975 ;
    RECT 53.975 14.665 54.245 14.735 ;
    RECT 53.975 15.425 54.245 15.495 ;
    RECT 53.975 16.185 54.245 16.255 ;
    RECT 53.975 16.945 54.245 17.015 ;
    RECT 53.975 17.705 54.245 17.775 ;
    RECT 53.975 18.465 54.245 18.535 ;
    RECT 53.975 19.225 54.245 19.295 ;
    RECT 53.975 19.985 54.245 20.055 ;
    RECT 53.975 20.745 54.245 20.815 ;
    RECT 53.975 21.505 54.245 21.575 ;
    RECT 53.975 22.265 54.245 22.335 ;
    RECT 53.975 23.025 54.245 23.095 ;
    RECT 56.07 11.625 56.34 11.695 ;
    RECT 56.07 12.385 56.34 12.455 ;
    RECT 56.07 13.145 56.34 13.215 ;
    RECT 56.07 13.905 56.34 13.975 ;
    RECT 56.07 14.665 56.34 14.735 ;
    RECT 56.07 15.425 56.34 15.495 ;
    RECT 56.07 16.185 56.34 16.255 ;
    RECT 56.07 16.945 56.34 17.015 ;
    RECT 56.07 17.705 56.34 17.775 ;
    RECT 56.07 18.465 56.34 18.535 ;
    RECT 56.07 19.225 56.34 19.295 ;
    RECT 56.07 19.985 56.34 20.055 ;
    RECT 56.07 20.745 56.34 20.815 ;
    RECT 56.07 21.505 56.34 21.575 ;
    RECT 56.07 22.265 56.34 22.335 ;
    RECT 56.07 23.025 56.34 23.095 ;
    RECT 79.54 11.625 79.61 11.695 ;
    RECT 79.54 12.385 79.61 12.455 ;
    RECT 79.54 13.145 79.61 13.215 ;
    RECT 79.54 13.905 79.61 13.975 ;
    RECT 79.54 14.665 79.61 14.735 ;
    RECT 79.54 15.425 79.61 15.495 ;
    RECT 79.54 16.185 79.61 16.255 ;
    RECT 79.54 16.945 79.61 17.015 ;
    RECT 79.54 17.705 79.61 17.775 ;
    RECT 79.54 18.465 79.61 18.535 ;
    RECT 79.54 19.225 79.61 19.295 ;
    RECT 79.54 19.985 79.61 20.055 ;
    RECT 79.54 20.745 79.61 20.815 ;
    RECT 79.54 21.505 79.61 21.575 ;
    RECT 79.54 22.265 79.61 22.335 ;
    RECT 79.54 23.025 79.61 23.095 ;
    RECT 80.525 11.625 80.595 11.695 ;
    RECT 80.525 12.385 80.595 12.455 ;
    RECT 80.525 13.145 80.595 13.215 ;
    RECT 80.525 13.905 80.595 13.975 ;
    RECT 80.525 14.665 80.595 14.735 ;
    RECT 80.525 15.425 80.785 15.495 ;
    RECT 80.525 16.185 80.595 16.255 ;
    RECT 80.525 16.945 80.595 17.015 ;
    RECT 80.525 17.705 80.595 17.775 ;
    RECT 80.525 18.465 80.595 18.535 ;
    RECT 80.525 19.225 80.595 19.295 ;
    RECT 80.525 19.985 80.595 20.055 ;
    RECT 80.525 20.745 80.595 20.815 ;
    RECT 80.525 21.505 80.595 21.575 ;
    RECT 80.525 22.265 80.595 22.335 ;
    RECT 80.525 23.025 80.595 23.095 ;
    RECT 80.715 11.625 80.785 11.695 ;
    RECT 80.715 12.385 80.785 12.455 ;
    RECT 80.715 13.145 80.785 13.215 ;
    RECT 80.715 13.905 80.785 13.975 ;
    RECT 80.715 14.665 80.785 14.735 ;
    RECT 80.715 16.185 80.785 16.255 ;
    RECT 80.715 16.945 80.785 17.015 ;
    RECT 80.715 17.705 80.785 17.775 ;
    RECT 80.715 18.465 80.785 18.535 ;
    RECT 80.715 19.225 80.785 19.295 ;
    RECT 80.715 19.985 80.785 20.055 ;
    RECT 80.715 20.745 80.785 20.815 ;
    RECT 80.715 21.505 80.785 21.575 ;
    RECT 80.715 22.265 80.785 22.335 ;
    RECT 80.715 23.025 80.785 23.095 ;
    RECT 48.415 11.005 48.625 11.075 ;
    RECT 45.62 11.005 45.83 11.075 ;
    RECT 44.225 11.005 44.435 11.075 ;
    RECT 42.825 11.005 43.035 11.075 ;
    RECT 40.03 11.005 40.24 11.075 ;
    RECT 38.635 11.005 38.845 11.075 ;
    RECT 37.24 11.005 37.45 11.075 ;
    RECT 33.045 11.005 33.255 11.075 ;
    RECT 31.65 11.005 31.86 11.075 ;
    RECT 28.855 11.005 29.065 11.075 ;
    RECT 27.455 11.005 27.665 11.075 ;
    RECT 74.97 109.98 75.18 110.05 ;
    RECT 73.57 109.98 73.78 110.05 ;
    RECT 70.77 109.98 70.98 110.05 ;
    RECT 69.37 109.98 69.58 110.05 ;
    RECT 67.975 109.98 68.185 110.05 ;
    RECT 63.785 109.98 63.995 110.05 ;
    RECT 62.385 110.155 62.595 110.365 ;
    RECT 58.195 109.98 58.405 110.05 ;
    RECT 56.8 109.98 57.01 110.05 ;
    RECT 53.305 109.98 53.515 110.05 ;
    RECT 51.91 109.98 52.12 110.05 ;
    RECT 30.67 108.125 30.74 108.195 ;
    RECT 50.93 108.125 51.0 108.195 ;
    RECT 53.975 108.125 54.245 108.195 ;
    RECT 56.07 108.125 56.34 108.195 ;
    RECT 79.575 108.125 79.645 108.195 ;
    RECT 30.67 107.365 30.74 107.435 ;
    RECT 50.93 107.365 51.0 107.435 ;
    RECT 53.975 107.365 54.245 107.435 ;
    RECT 56.07 107.365 56.34 107.435 ;
    RECT 79.575 107.365 79.645 107.435 ;
    RECT 30.67 106.605 30.74 106.675 ;
    RECT 50.93 106.605 51.0 106.675 ;
    RECT 53.975 106.605 54.245 106.675 ;
    RECT 56.07 106.605 56.34 106.675 ;
    RECT 79.575 106.605 79.645 106.675 ;
    RECT 30.67 105.845 30.74 105.915 ;
    RECT 50.93 105.845 51.0 105.915 ;
    RECT 53.975 105.845 54.245 105.915 ;
    RECT 56.07 105.845 56.34 105.915 ;
    RECT 79.575 105.845 79.645 105.915 ;
    RECT 30.67 105.085 30.74 105.155 ;
    RECT 50.93 105.085 51.0 105.155 ;
    RECT 53.975 105.085 54.245 105.155 ;
    RECT 56.07 105.085 56.34 105.155 ;
    RECT 79.575 105.085 79.645 105.155 ;
    RECT 30.67 104.325 30.74 104.395 ;
    RECT 50.93 104.325 51.0 104.395 ;
    RECT 53.975 104.325 54.245 104.395 ;
    RECT 56.07 104.325 56.34 104.395 ;
    RECT 79.575 104.325 79.645 104.395 ;
    RECT 30.67 103.565 30.74 103.635 ;
    RECT 50.93 103.565 51.0 103.635 ;
    RECT 53.975 103.565 54.245 103.635 ;
    RECT 56.07 103.565 56.34 103.635 ;
    RECT 79.575 103.565 79.645 103.635 ;
    RECT 30.67 102.805 30.74 102.875 ;
    RECT 50.93 102.805 51.0 102.875 ;
    RECT 53.975 102.805 54.245 102.875 ;
    RECT 56.07 102.805 56.34 102.875 ;
    RECT 79.575 102.805 79.645 102.875 ;
    RECT 30.67 102.045 30.74 102.115 ;
    RECT 50.93 102.045 51.0 102.115 ;
    RECT 53.975 102.045 54.245 102.115 ;
    RECT 56.07 102.045 56.34 102.115 ;
    RECT 79.575 102.045 79.645 102.115 ;
    RECT 30.67 101.285 30.74 101.355 ;
    RECT 50.93 101.285 51.0 101.355 ;
    RECT 53.975 101.285 54.245 101.355 ;
    RECT 56.07 101.285 56.34 101.355 ;
    RECT 79.575 101.285 79.645 101.355 ;
    RECT 30.67 100.525 30.74 100.595 ;
    RECT 50.93 100.525 51.0 100.595 ;
    RECT 53.975 100.525 54.245 100.595 ;
    RECT 56.07 100.525 56.34 100.595 ;
    RECT 79.575 100.525 79.645 100.595 ;
    RECT 30.67 99.765 30.74 99.835 ;
    RECT 50.93 99.765 51.0 99.835 ;
    RECT 53.975 99.765 54.245 99.835 ;
    RECT 56.07 99.765 56.34 99.835 ;
    RECT 79.575 99.765 79.645 99.835 ;
    RECT 30.67 99.005 30.74 99.075 ;
    RECT 50.93 99.005 51.0 99.075 ;
    RECT 53.975 99.005 54.245 99.075 ;
    RECT 56.07 99.005 56.34 99.075 ;
    RECT 79.575 99.005 79.645 99.075 ;
    RECT 30.67 98.245 30.74 98.315 ;
    RECT 50.93 98.245 51.0 98.315 ;
    RECT 53.975 98.245 54.245 98.315 ;
    RECT 56.07 98.245 56.34 98.315 ;
    RECT 79.575 98.245 79.645 98.315 ;
    RECT 30.67 97.485 30.74 97.555 ;
    RECT 50.93 97.485 51.0 97.555 ;
    RECT 53.975 97.485 54.245 97.555 ;
    RECT 56.07 97.485 56.34 97.555 ;
    RECT 79.575 97.485 79.645 97.555 ;
    RECT 30.67 96.725 30.74 96.795 ;
    RECT 50.93 96.725 51.0 96.795 ;
    RECT 53.975 96.725 54.245 96.795 ;
    RECT 56.07 96.725 56.34 96.795 ;
    RECT 79.575 96.725 79.645 96.795 ;
    RECT 30.67 95.965 30.74 96.035 ;
    RECT 50.93 95.965 51.0 96.035 ;
    RECT 53.975 95.965 54.245 96.035 ;
    RECT 56.07 95.965 56.34 96.035 ;
    RECT 79.575 95.965 79.645 96.035 ;
    RECT 30.67 95.205 30.74 95.275 ;
    RECT 50.93 95.205 51.0 95.275 ;
    RECT 53.975 95.205 54.245 95.275 ;
    RECT 56.07 95.205 56.34 95.275 ;
    RECT 79.575 95.205 79.645 95.275 ;
    RECT 30.67 94.445 30.74 94.515 ;
    RECT 50.93 94.445 51.0 94.515 ;
    RECT 53.975 94.445 54.245 94.515 ;
    RECT 56.07 94.445 56.34 94.515 ;
    RECT 79.575 94.445 79.645 94.515 ;
    RECT 30.67 93.685 30.74 93.755 ;
    RECT 50.93 93.685 51.0 93.755 ;
    RECT 53.975 93.685 54.245 93.755 ;
    RECT 56.07 93.685 56.34 93.755 ;
    RECT 79.575 93.685 79.645 93.755 ;
    RECT 30.67 92.925 30.74 92.995 ;
    RECT 50.93 92.925 51.0 92.995 ;
    RECT 53.975 92.925 54.245 92.995 ;
    RECT 56.07 92.925 56.34 92.995 ;
    RECT 79.575 92.925 79.645 92.995 ;
    RECT 30.67 92.165 30.74 92.235 ;
    RECT 50.93 92.165 51.0 92.235 ;
    RECT 53.975 92.165 54.245 92.235 ;
    RECT 56.07 92.165 56.34 92.235 ;
    RECT 79.575 92.165 79.645 92.235 ;
    RECT 30.67 91.405 30.74 91.475 ;
    RECT 50.93 91.405 51.0 91.475 ;
    RECT 53.975 91.405 54.245 91.475 ;
    RECT 56.07 91.405 56.34 91.475 ;
    RECT 79.575 91.405 79.645 91.475 ;
    RECT 30.67 90.645 30.74 90.715 ;
    RECT 50.93 90.645 51.0 90.715 ;
    RECT 53.975 90.645 54.245 90.715 ;
    RECT 56.07 90.645 56.34 90.715 ;
    RECT 79.575 90.645 79.645 90.715 ;
    RECT 30.67 89.885 30.74 89.955 ;
    RECT 50.93 89.885 51.0 89.955 ;
    RECT 53.975 89.885 54.245 89.955 ;
    RECT 56.07 89.885 56.34 89.955 ;
    RECT 79.575 89.885 79.645 89.955 ;
    RECT 30.67 89.125 30.74 89.195 ;
    RECT 50.93 89.125 51.0 89.195 ;
    RECT 53.975 89.125 54.245 89.195 ;
    RECT 56.07 89.125 56.34 89.195 ;
    RECT 79.575 89.125 79.645 89.195 ;
    RECT 30.67 88.365 30.74 88.435 ;
    RECT 50.93 88.365 51.0 88.435 ;
    RECT 53.975 88.365 54.245 88.435 ;
    RECT 56.07 88.365 56.34 88.435 ;
    RECT 79.575 88.365 79.645 88.435 ;
    RECT 30.67 87.605 30.74 87.675 ;
    RECT 50.93 87.605 51.0 87.675 ;
    RECT 53.975 87.605 54.245 87.675 ;
    RECT 56.07 87.605 56.34 87.675 ;
    RECT 79.575 87.605 79.645 87.675 ;
    RECT 30.67 108.885 30.74 108.955 ;
    RECT 50.93 108.885 51.0 108.955 ;
    RECT 53.975 108.885 54.245 108.955 ;
    RECT 56.07 108.885 56.34 108.955 ;
    RECT 79.575 108.885 79.645 108.955 ;
    RECT 82.65 60.415 82.86 60.485 ;
    RECT 81.25 60.415 81.46 60.485 ;
    RECT 78.455 60.415 78.665 60.485 ;
    RECT 77.055 60.415 77.265 60.485 ;
    RECT 75.67 60.555 75.88 60.625 ;
    RECT 75.67 59.955 75.88 60.025 ;
    RECT 72.87 60.415 73.08 60.485 ;
    RECT 71.47 60.415 71.68 60.485 ;
    RECT 70.07 60.415 70.28 60.485 ;
    RECT 67.275 60.415 67.485 60.485 ;
    RECT 65.88 60.415 66.09 60.485 ;
    RECT 64.48 60.415 64.69 60.485 ;
    RECT 61.69 60.415 61.9 60.485 ;
    RECT 60.295 60.415 60.505 60.485 ;
    RECT 47.715 110.155 47.925 110.365 ;
    RECT 46.32 109.98 46.53 110.05 ;
    RECT 42.13 109.98 42.34 110.05 ;
    RECT 40.73 109.98 40.94 110.05 ;
    RECT 39.335 109.98 39.545 110.05 ;
    RECT 36.54 109.98 36.75 110.05 ;
    RECT 35.14 109.98 35.35 110.05 ;
    RECT 82.65 109.505 82.86 109.575 ;
    RECT 81.25 109.485 81.46 109.555 ;
    RECT 78.455 109.485 78.665 109.555 ;
    RECT 77.055 109.485 77.265 109.555 ;
    RECT 75.67 109.335 75.88 109.405 ;
    RECT 72.87 109.485 73.08 109.555 ;
    RECT 71.47 109.485 71.68 109.555 ;
    RECT 70.07 109.485 70.28 109.555 ;
    RECT 67.275 109.485 67.485 109.555 ;
    RECT 65.88 109.485 66.09 109.555 ;
    RECT 64.48 109.485 64.69 109.555 ;
    RECT 61.69 109.485 61.9 109.555 ;
    RECT 60.295 109.485 60.505 109.555 ;
    RECT 56.1 109.485 56.31 109.555 ;
    RECT 54.005 109.485 54.215 109.555 ;
    RECT 49.815 109.485 50.025 109.555 ;
    RECT 48.415 109.485 48.625 109.555 ;
    RECT 45.62 109.485 45.83 109.555 ;
    RECT 44.225 109.485 44.435 109.555 ;
    RECT 42.825 109.485 43.035 109.555 ;
    RECT 40.03 109.485 40.24 109.555 ;
    RECT 38.635 109.485 38.845 109.555 ;
    RECT 37.24 109.485 37.45 109.555 ;
    RECT 34.445 109.335 34.655 109.405 ;
    RECT 33.045 109.485 33.255 109.555 ;
    RECT 31.65 109.485 31.86 109.555 ;
    RECT 28.855 109.485 29.065 109.555 ;
    RECT 27.455 109.485 27.665 109.555 ;
    RECT 77.755 109.655 77.965 109.725 ;
    RECT 76.36 109.655 76.57 109.725 ;
    RECT 72.17 109.655 72.38 109.725 ;
    RECT 66.58 109.655 66.79 109.725 ;
    RECT 65.18 109.655 65.39 109.725 ;
    RECT 60.99 109.655 61.2 109.725 ;
    RECT 55.4 109.655 55.61 109.725 ;
    RECT 54.705 109.655 54.915 109.725 ;
    RECT 49.115 109.655 49.325 109.725 ;
    RECT 44.925 109.655 45.135 109.725 ;
    RECT 43.525 109.655 43.735 109.725 ;
    RECT 37.935 109.655 38.145 109.725 ;
    RECT 33.745 109.655 33.955 109.725 ;
    RECT 32.345 109.655 32.555 109.725 ;
    RECT 77.755 60.12 77.965 60.19 ;
    RECT 76.36 60.12 76.57 60.19 ;
    RECT 72.17 60.12 72.38 60.19 ;
    RECT 66.58 60.12 66.79 60.19 ;
    RECT 65.18 60.12 65.39 60.19 ;
    RECT 60.99 60.12 61.2 60.19 ;
    RECT 55.4 60.12 55.61 60.19 ;
    RECT 54.705 60.12 54.915 60.19 ;
    RECT 49.115 60.12 49.325 60.19 ;
    RECT 44.925 60.12 45.135 60.19 ;
    RECT 32.345 110.485 32.555 110.695 ;
    RECT 26.915 10.055 27.125 10.265 ;
    RECT 83.09 10.055 83.3 10.265 ;
    RECT 77.755 10.055 77.965 10.265 ;
    RECT 76.36 10.055 76.57 10.265 ;
    RECT 72.17 10.055 72.38 10.265 ;
    RECT 66.58 10.055 66.79 10.265 ;
    RECT 65.18 10.055 65.39 10.265 ;
    RECT 60.99 10.055 61.2 10.265 ;
    RECT 55.4 10.055 55.61 10.265 ;
    RECT 54.705 10.055 54.915 10.265 ;
    RECT 49.115 10.055 49.325 10.265 ;
    RECT 44.925 10.055 45.135 10.265 ;
    RECT 43.525 10.055 43.735 10.265 ;
    RECT 37.935 10.055 38.145 10.265 ;
    RECT 33.745 10.055 33.955 10.265 ;
    RECT 32.345 10.055 32.555 10.265 ;
    RECT 58.895 10.055 59.105 10.265 ;
    RECT 80.55 10.055 80.76 10.265 ;
    RECT 51.21 10.055 51.42 10.265 ;
    RECT 29.555 10.055 29.765 10.265 ;
    RECT 78.455 11.175 78.665 11.245 ;
    RECT 77.055 11.175 77.265 11.245 ;
    RECT 72.87 11.175 73.08 11.245 ;
    RECT 71.47 11.175 71.68 11.245 ;
    RECT 70.07 11.175 70.28 11.245 ;
    RECT 67.275 11.175 67.485 11.245 ;
    RECT 65.88 11.175 66.09 11.245 ;
    RECT 64.48 11.175 64.69 11.245 ;
    RECT 61.69 11.175 61.9 11.245 ;
    RECT 60.295 11.175 60.505 11.245 ;
    RECT 56.1 11.175 56.31 11.245 ;
    RECT 54.005 11.175 54.215 11.245 ;
    RECT 49.815 11.175 50.025 11.245 ;
    RECT 48.415 11.175 48.625 11.245 ;
    RECT 45.62 11.175 45.83 11.245 ;
    RECT 44.225 11.175 44.435 11.245 ;
    RECT 42.825 11.175 43.035 11.245 ;
    RECT 40.03 11.175 40.24 11.245 ;
    RECT 38.635 11.175 38.845 11.245 ;
    RECT 37.24 11.175 37.45 11.245 ;
    RECT 56.1 60.415 56.31 60.485 ;
    RECT 54.005 60.415 54.215 60.485 ;
    RECT 49.815 60.415 50.025 60.485 ;
    RECT 33.045 11.175 33.255 11.245 ;
    RECT 48.415 60.415 48.625 60.485 ;
    RECT 45.62 60.415 45.83 60.485 ;
    RECT 31.65 11.175 31.86 11.245 ;
    RECT 44.225 60.415 44.435 60.485 ;
    RECT 42.825 60.415 43.035 60.485 ;
    RECT 40.03 60.415 40.24 60.485 ;
    RECT 38.635 60.415 38.845 60.485 ;
    RECT 37.24 60.415 37.45 60.485 ;
    RECT 34.445 60.555 34.655 60.625 ;
    RECT 34.445 59.955 34.655 60.025 ;
    RECT 33.045 60.415 33.255 60.485 ;
    RECT 31.65 60.415 31.86 60.485 ;
    RECT 28.855 60.415 29.065 60.485 ;
    RECT 27.455 60.415 27.665 60.485 ;
    RECT 77.755 60.275 77.965 60.345 ;
    RECT 76.36 60.275 76.57 60.345 ;
    RECT 72.17 60.275 72.38 60.345 ;
    RECT 66.58 60.275 66.79 60.345 ;
    RECT 65.18 60.275 65.39 60.345 ;
    RECT 60.99 60.275 61.2 60.345 ;
    RECT 55.4 60.275 55.61 60.345 ;
    RECT 54.705 60.275 54.915 60.345 ;
    RECT 49.115 60.275 49.325 60.345 ;
    RECT 44.925 60.275 45.135 60.345 ;
    RECT 43.525 60.275 43.735 60.345 ;
    RECT 37.935 60.275 38.145 60.345 ;
    RECT 33.745 60.275 33.955 60.345 ;
    RECT 32.345 60.275 32.555 60.345 ;
    RECT 77.755 10.752 77.965 10.822 ;
    RECT 76.36 10.752 76.57 10.822 ;
    RECT 72.17 10.752 72.38 10.822 ;
    RECT 66.58 10.752 66.79 10.822 ;
    RECT 65.18 10.752 65.39 10.822 ;
    RECT 60.99 10.752 61.2 10.822 ;
    RECT 55.4 10.752 55.61 10.822 ;
    RECT 54.705 10.752 54.915 10.822 ;
    RECT 49.115 10.752 49.325 10.822 ;
    RECT 44.925 10.752 45.135 10.822 ;
    RECT 43.525 10.752 43.735 10.822 ;
    RECT 37.935 10.752 38.145 10.822 ;
    RECT 33.745 10.752 33.955 10.822 ;
    RECT 32.345 10.752 32.555 10.822 ;
    RECT 43.525 60.12 43.735 60.19 ;
    RECT 37.935 60.12 38.145 60.19 ;
    RECT 33.745 60.12 33.955 60.19 ;
    RECT 32.345 60.12 32.555 60.19 ;
    RECT 79.855 60.555 80.065 60.625 ;
    RECT 79.855 59.955 80.065 60.025 ;
    RECT 74.27 60.555 74.48 60.625 ;
    RECT 74.27 59.955 74.48 60.025 ;
    RECT 68.675 59.955 68.885 60.025 ;
    RECT 63.085 60.555 63.295 60.625 ;
    RECT 63.085 59.955 63.295 60.025 ;
    RECT 57.5 60.555 57.71 60.625 ;
    RECT 57.5 59.955 57.71 60.025 ;
    RECT 52.61 60.555 52.82 60.625 ;
    RECT 52.61 59.955 52.82 60.025 ;
    RECT 47.02 60.555 47.23 60.625 ;
    RECT 47.02 59.955 47.23 60.025 ;
    RECT 41.43 59.955 41.64 60.025 ;
    RECT 35.84 60.555 36.05 60.625 ;
    RECT 35.84 59.955 36.05 60.025 ;
    RECT 30.25 60.555 30.46 60.625 ;
    RECT 30.25 59.955 30.46 60.025 ;
    RECT 79.855 109.335 80.065 109.405 ;
    RECT 74.27 109.335 74.48 109.405 ;
    RECT 68.675 109.335 68.885 109.405 ;
    RECT 63.085 109.335 63.295 109.405 ;
    RECT 57.5 109.335 57.71 109.405 ;
    RECT 52.61 109.335 52.82 109.405 ;
    RECT 47.02 109.335 47.23 109.405 ;
    RECT 41.43 109.335 41.64 109.405 ;
    RECT 35.84 109.335 36.05 109.405 ;
    RECT 30.25 109.335 30.46 109.405 ;
    RECT 77.755 110.485 77.965 110.695 ;
    RECT 76.36 110.485 76.57 110.695 ;
    RECT 72.17 110.485 72.38 110.695 ;
    RECT 66.58 110.485 66.79 110.695 ;
    RECT 65.18 110.485 65.39 110.695 ;
    RECT 60.99 110.485 61.2 110.695 ;
    RECT 55.4 110.485 55.61 110.695 ;
    RECT 54.705 110.485 54.915 110.695 ;
    RECT 49.115 110.485 49.325 110.695 ;
    RECT 44.925 110.485 45.135 110.695 ;
    RECT 43.525 110.485 43.735 110.695 ;
    RECT 37.935 110.485 38.145 110.695 ;
    RECT 33.745 110.485 33.955 110.695 ;
    RECT 30.67 86.845 30.74 86.915 ;
    RECT 50.93 86.845 51.0 86.915 ;
    RECT 53.975 86.845 54.245 86.915 ;
    RECT 56.07 86.845 56.34 86.915 ;
    RECT 79.575 86.845 79.645 86.915 ;
    RECT 30.67 86.085 30.74 86.155 ;
    RECT 50.93 86.085 51.0 86.155 ;
    RECT 53.975 86.085 54.245 86.155 ;
    RECT 56.07 86.085 56.34 86.155 ;
    RECT 79.575 86.085 79.645 86.155 ;
    RECT 30.67 85.325 30.74 85.395 ;
    RECT 50.93 85.325 51.0 85.395 ;
    RECT 53.975 85.325 54.245 85.395 ;
    RECT 56.07 85.325 56.34 85.395 ;
    RECT 79.575 85.325 79.645 85.395 ;
    RECT 30.67 84.565 30.74 84.635 ;
    RECT 50.93 84.565 51.0 84.635 ;
    RECT 53.975 84.565 54.245 84.635 ;
    RECT 56.07 84.565 56.34 84.635 ;
    RECT 79.575 84.565 79.645 84.635 ;
    RECT 30.67 83.805 30.74 83.875 ;
    RECT 50.93 83.805 51.0 83.875 ;
    RECT 53.975 83.805 54.245 83.875 ;
    RECT 56.07 83.805 56.34 83.875 ;
    RECT 79.575 83.805 79.645 83.875 ;
    RECT 30.67 83.045 30.74 83.115 ;
    RECT 50.93 83.045 51.0 83.115 ;
    RECT 53.975 83.045 54.245 83.115 ;
    RECT 56.07 83.045 56.34 83.115 ;
    RECT 79.575 83.045 79.645 83.115 ;
    RECT 30.67 82.285 30.74 82.355 ;
    RECT 50.93 82.285 51.0 82.355 ;
    RECT 53.975 82.285 54.245 82.355 ;
    RECT 56.07 82.285 56.34 82.355 ;
    RECT 79.575 82.285 79.645 82.355 ;
    RECT 30.67 81.525 30.74 81.595 ;
    RECT 50.93 81.525 51.0 81.595 ;
    RECT 53.975 81.525 54.245 81.595 ;
    RECT 56.07 81.525 56.34 81.595 ;
    RECT 79.575 81.525 79.645 81.595 ;
    RECT 30.67 80.765 30.74 80.835 ;
    RECT 50.93 80.765 51.0 80.835 ;
    RECT 53.975 80.765 54.245 80.835 ;
    RECT 56.07 80.765 56.34 80.835 ;
    RECT 79.575 80.765 79.645 80.835 ;
    RECT 30.67 80.005 30.74 80.075 ;
    RECT 50.93 80.005 51.0 80.075 ;
    RECT 53.975 80.005 54.245 80.075 ;
    RECT 56.07 80.005 56.34 80.075 ;
    RECT 79.575 80.005 79.645 80.075 ;
    RECT 30.67 79.245 30.74 79.315 ;
    RECT 50.93 79.245 51.0 79.315 ;
    RECT 53.975 79.245 54.245 79.315 ;
    RECT 56.07 79.245 56.34 79.315 ;
    RECT 79.575 79.245 79.645 79.315 ;
    RECT 30.67 78.485 30.74 78.555 ;
    RECT 50.93 78.485 51.0 78.555 ;
    RECT 53.975 78.485 54.245 78.555 ;
    RECT 56.07 78.485 56.34 78.555 ;
    RECT 79.575 78.485 79.645 78.555 ;
    RECT 30.67 77.725 30.74 77.795 ;
    RECT 50.93 77.725 51.0 77.795 ;
    RECT 53.975 77.725 54.245 77.795 ;
    RECT 56.07 77.725 56.34 77.795 ;
    RECT 79.575 77.725 79.645 77.795 ;
    RECT 30.67 76.965 30.74 77.035 ;
    RECT 50.93 76.965 51.0 77.035 ;
    RECT 53.975 76.965 54.245 77.035 ;
    RECT 56.07 76.965 56.34 77.035 ;
    RECT 79.575 76.965 79.645 77.035 ;
    RECT 30.67 76.205 30.74 76.275 ;
    RECT 50.93 76.205 51.0 76.275 ;
    RECT 53.975 76.205 54.245 76.275 ;
    RECT 56.07 76.205 56.34 76.275 ;
    RECT 79.575 76.205 79.645 76.275 ;
    RECT 30.67 75.445 30.74 75.515 ;
    RECT 50.93 75.445 51.0 75.515 ;
    RECT 53.975 75.445 54.245 75.515 ;
    RECT 56.07 75.445 56.34 75.515 ;
    RECT 79.575 75.445 79.645 75.515 ;
    RECT 30.67 74.685 30.74 74.755 ;
    RECT 50.93 74.685 51.0 74.755 ;
    RECT 53.975 74.685 54.245 74.755 ;
    RECT 56.07 74.685 56.34 74.755 ;
    RECT 79.575 74.685 79.645 74.755 ;
    RECT 30.67 73.925 30.74 73.995 ;
    RECT 50.93 73.925 51.0 73.995 ;
    RECT 53.975 73.925 54.245 73.995 ;
    RECT 56.07 73.925 56.34 73.995 ;
    RECT 79.575 73.925 79.645 73.995 ;
    RECT 30.67 73.165 30.74 73.235 ;
    RECT 50.93 73.165 51.0 73.235 ;
    RECT 53.975 73.165 54.245 73.235 ;
    RECT 56.07 73.165 56.34 73.235 ;
    RECT 79.575 73.165 79.645 73.235 ;
    RECT 30.67 72.405 30.74 72.475 ;
    RECT 50.93 72.405 51.0 72.475 ;
    RECT 53.975 72.405 54.245 72.475 ;
    RECT 56.07 72.405 56.34 72.475 ;
    RECT 79.575 72.405 79.645 72.475 ;
    RECT 30.67 71.645 30.74 71.715 ;
    RECT 50.93 71.645 51.0 71.715 ;
    RECT 53.975 71.645 54.245 71.715 ;
    RECT 56.07 71.645 56.34 71.715 ;
    RECT 79.575 71.645 79.645 71.715 ;
    RECT 30.67 70.885 30.74 70.955 ;
    RECT 50.93 70.885 51.0 70.955 ;
    RECT 53.975 70.885 54.245 70.955 ;
    RECT 56.07 70.885 56.34 70.955 ;
    RECT 79.575 70.885 79.645 70.955 ;
    RECT 30.67 70.125 30.74 70.195 ;
    RECT 50.93 70.125 51.0 70.195 ;
    RECT 53.975 70.125 54.245 70.195 ;
    RECT 56.07 70.125 56.34 70.195 ;
    RECT 79.575 70.125 79.645 70.195 ;
    RECT 30.67 69.365 30.74 69.435 ;
    RECT 50.93 69.365 51.0 69.435 ;
    RECT 53.975 69.365 54.245 69.435 ;
    RECT 56.07 69.365 56.34 69.435 ;
    RECT 79.575 69.365 79.645 69.435 ;
    RECT 30.67 68.605 30.74 68.675 ;
    RECT 50.93 68.605 51.0 68.675 ;
    RECT 53.975 68.605 54.245 68.675 ;
    RECT 56.07 68.605 56.34 68.675 ;
    RECT 79.575 68.605 79.645 68.675 ;
    RECT 30.67 67.845 30.74 67.915 ;
    RECT 50.93 67.845 51.0 67.915 ;
    RECT 53.975 67.845 54.245 67.915 ;
    RECT 56.07 67.845 56.34 67.915 ;
    RECT 79.575 67.845 79.645 67.915 ;
    RECT 30.67 67.085 30.74 67.155 ;
    RECT 50.93 67.085 51.0 67.155 ;
    RECT 53.975 67.085 54.245 67.155 ;
    RECT 56.07 67.085 56.34 67.155 ;
    RECT 79.575 67.085 79.645 67.155 ;
    RECT 30.67 66.325 30.74 66.395 ;
    RECT 50.93 66.325 51.0 66.395 ;
    RECT 53.975 66.325 54.245 66.395 ;
    RECT 56.07 66.325 56.34 66.395 ;
    RECT 79.575 66.325 79.645 66.395 ;
    RECT 30.67 65.565 30.74 65.635 ;
    RECT 50.93 65.565 51.0 65.635 ;
    RECT 53.975 65.565 54.245 65.635 ;
    RECT 56.07 65.565 56.34 65.635 ;
    RECT 79.575 65.565 79.645 65.635 ;
    RECT 30.67 64.805 30.74 64.875 ;
    RECT 50.93 64.805 51.0 64.875 ;
    RECT 53.975 64.805 54.245 64.875 ;
    RECT 56.07 64.805 56.34 64.875 ;
    RECT 79.575 64.805 79.645 64.875 ;
    RECT 30.67 64.045 30.74 64.115 ;
    RECT 50.93 64.045 51.0 64.115 ;
    RECT 53.975 64.045 54.245 64.115 ;
    RECT 56.07 64.045 56.34 64.115 ;
    RECT 79.575 64.045 79.645 64.115 ;
    RECT 30.67 63.285 30.74 63.355 ;
    RECT 50.93 63.285 51.0 63.355 ;
    RECT 53.975 63.285 54.245 63.355 ;
    RECT 56.07 63.285 56.34 63.355 ;
    RECT 79.575 63.285 79.645 63.355 ;
    RECT 30.67 62.525 30.74 62.595 ;
    RECT 50.93 62.525 51.0 62.595 ;
    RECT 53.975 62.525 54.245 62.595 ;
    RECT 56.07 62.525 56.34 62.595 ;
    RECT 79.575 62.525 79.645 62.595 ;
    RECT 30.67 61.765 30.74 61.835 ;
    RECT 50.93 61.765 51.0 61.835 ;
    RECT 53.975 61.765 54.245 61.835 ;
    RECT 56.07 61.765 56.34 61.835 ;
    RECT 79.575 61.765 79.645 61.835 ;
    RECT 30.67 61.005 30.74 61.075 ;
    RECT 50.93 61.005 51.0 61.075 ;
    RECT 53.975 61.005 54.245 61.075 ;
    RECT 56.07 61.005 56.34 61.075 ;
    RECT 79.575 61.005 79.645 61.075 ;
    RECT 42.095 60.555 42.365 60.625 ;
    RECT 67.945 60.555 68.215 60.625 ;
    RECT 30.67 59.505 30.74 59.575 ;
    RECT 50.93 59.505 51.0 59.575 ;
    RECT 53.975 59.505 54.245 59.575 ;
    RECT 56.07 59.505 56.34 59.575 ;
    RECT 79.575 59.505 79.645 59.575 ;
    RECT 30.67 58.745 30.74 58.815 ;
    RECT 50.93 58.745 51.0 58.815 ;
    RECT 53.975 58.745 54.245 58.815 ;
    RECT 56.07 58.745 56.34 58.815 ;
    RECT 79.575 58.745 79.645 58.815 ;
    RECT 30.67 57.985 30.74 58.055 ;
    RECT 50.93 57.985 51.0 58.055 ;
    RECT 53.975 57.985 54.245 58.055 ;
    RECT 56.07 57.985 56.34 58.055 ;
    RECT 79.575 57.985 79.645 58.055 ;
    RECT 30.67 57.225 30.74 57.295 ;
    RECT 50.93 57.225 51.0 57.295 ;
    RECT 53.975 57.225 54.245 57.295 ;
    RECT 56.07 57.225 56.34 57.295 ;
    RECT 79.575 57.225 79.645 57.295 ;
    RECT 30.67 56.465 30.74 56.535 ;
    RECT 50.93 56.465 51.0 56.535 ;
    RECT 53.975 56.465 54.245 56.535 ;
    RECT 56.07 56.465 56.34 56.535 ;
    RECT 79.575 56.465 79.645 56.535 ;
    RECT 30.67 55.705 30.74 55.775 ;
    RECT 50.93 55.705 51.0 55.775 ;
    RECT 53.975 55.705 54.245 55.775 ;
    RECT 56.07 55.705 56.34 55.775 ;
    RECT 79.575 55.705 79.645 55.775 ;
    RECT 30.67 54.945 30.74 55.015 ;
    RECT 50.93 54.945 51.0 55.015 ;
    RECT 53.975 54.945 54.245 55.015 ;
    RECT 56.07 54.945 56.34 55.015 ;
    RECT 79.575 54.945 79.645 55.015 ;
    RECT 30.67 54.185 30.74 54.255 ;
    RECT 50.93 54.185 51.0 54.255 ;
    RECT 53.975 54.185 54.245 54.255 ;
    RECT 56.07 54.185 56.34 54.255 ;
    RECT 79.575 54.185 79.645 54.255 ;
    RECT 30.67 53.425 30.74 53.495 ;
    RECT 50.93 53.425 51.0 53.495 ;
    RECT 53.975 53.425 54.245 53.495 ;
    RECT 56.07 53.425 56.34 53.495 ;
    RECT 79.575 53.425 79.645 53.495 ;
    RECT 30.67 52.665 30.74 52.735 ;
    RECT 50.93 52.665 51.0 52.735 ;
    RECT 53.975 52.665 54.245 52.735 ;
    RECT 56.07 52.665 56.34 52.735 ;
    RECT 79.575 52.665 79.645 52.735 ;
    RECT 30.67 51.905 30.74 51.975 ;
    RECT 50.93 51.905 51.0 51.975 ;
    RECT 53.975 51.905 54.245 51.975 ;
    RECT 56.07 51.905 56.34 51.975 ;
    RECT 79.575 51.905 79.645 51.975 ;
    RECT 30.67 51.145 30.74 51.215 ;
    RECT 50.93 51.145 51.0 51.215 ;
    RECT 53.975 51.145 54.245 51.215 ;
    RECT 56.07 51.145 56.34 51.215 ;
    RECT 79.575 51.145 79.645 51.215 ;
    RECT 30.67 50.385 30.74 50.455 ;
    RECT 50.93 50.385 51.0 50.455 ;
    RECT 53.975 50.385 54.245 50.455 ;
    RECT 56.07 50.385 56.34 50.455 ;
    RECT 79.575 50.385 79.645 50.455 ;
    RECT 30.67 49.625 30.74 49.695 ;
    RECT 50.93 49.625 51.0 49.695 ;
    RECT 53.975 49.625 54.245 49.695 ;
    RECT 56.07 49.625 56.34 49.695 ;
    RECT 79.575 49.625 79.645 49.695 ;
    RECT 30.67 48.865 30.74 48.935 ;
    RECT 50.93 48.865 51.0 48.935 ;
    RECT 53.975 48.865 54.245 48.935 ;
    RECT 56.07 48.865 56.34 48.935 ;
    RECT 79.575 48.865 79.645 48.935 ;
    RECT 30.67 48.105 30.74 48.175 ;
    RECT 50.93 48.105 51.0 48.175 ;
    RECT 53.975 48.105 54.245 48.175 ;
    RECT 56.07 48.105 56.34 48.175 ;
    RECT 79.575 48.105 79.645 48.175 ;
    RECT 30.67 47.345 30.74 47.415 ;
    RECT 50.93 47.345 51.0 47.415 ;
    RECT 53.975 47.345 54.245 47.415 ;
    RECT 56.07 47.345 56.34 47.415 ;
    RECT 79.575 47.345 79.645 47.415 ;
    RECT 30.67 46.585 30.74 46.655 ;
    RECT 50.93 46.585 51.0 46.655 ;
    RECT 53.975 46.585 54.245 46.655 ;
    RECT 56.07 46.585 56.34 46.655 ;
    RECT 79.575 46.585 79.645 46.655 ;
    RECT 30.67 45.825 30.74 45.895 ;
    RECT 50.93 45.825 51.0 45.895 ;
    RECT 53.975 45.825 54.245 45.895 ;
    RECT 56.07 45.825 56.34 45.895 ;
    RECT 79.575 45.825 79.645 45.895 ;
    RECT 30.67 45.065 30.74 45.135 ;
    RECT 50.93 45.065 51.0 45.135 ;
    RECT 53.975 45.065 54.245 45.135 ;
    RECT 56.07 45.065 56.34 45.135 ;
    RECT 79.575 45.065 79.645 45.135 ;
    RECT 30.67 44.305 30.74 44.375 ;
    RECT 50.93 44.305 51.0 44.375 ;
    RECT 53.975 44.305 54.245 44.375 ;
    RECT 56.07 44.305 56.34 44.375 ;
    RECT 79.575 44.305 79.645 44.375 ;
    RECT 30.67 43.545 30.74 43.615 ;
    RECT 50.93 43.545 51.0 43.615 ;
    RECT 53.975 43.545 54.245 43.615 ;
    RECT 56.07 43.545 56.34 43.615 ;
    RECT 79.575 43.545 79.645 43.615 ;
    RECT 30.67 42.785 30.74 42.855 ;
    RECT 50.93 42.785 51.0 42.855 ;
    RECT 53.975 42.785 54.245 42.855 ;
    RECT 56.07 42.785 56.34 42.855 ;
    RECT 79.575 42.785 79.645 42.855 ;
    RECT 30.67 42.025 30.74 42.095 ;
    RECT 50.93 42.025 51.0 42.095 ;
    RECT 53.975 42.025 54.245 42.095 ;
    RECT 56.07 42.025 56.34 42.095 ;
    RECT 79.575 42.025 79.645 42.095 ;
    RECT 30.67 41.265 30.74 41.335 ;
    RECT 50.93 41.265 51.0 41.335 ;
    RECT 53.975 41.265 54.245 41.335 ;
    RECT 56.07 41.265 56.34 41.335 ;
    RECT 79.575 41.265 79.645 41.335 ;
    RECT 30.67 40.505 30.74 40.575 ;
    RECT 50.93 40.505 51.0 40.575 ;
    RECT 53.975 40.505 54.245 40.575 ;
    RECT 56.07 40.505 56.34 40.575 ;
    RECT 79.575 40.505 79.645 40.575 ;
    RECT 30.67 39.745 30.74 39.815 ;
    RECT 50.93 39.745 51.0 39.815 ;
    RECT 53.975 39.745 54.245 39.815 ;
    RECT 56.07 39.745 56.34 39.815 ;
    RECT 79.575 39.745 79.645 39.815 ;
    RECT 30.67 38.985 30.74 39.055 ;
    RECT 50.93 38.985 51.0 39.055 ;
    RECT 53.975 38.985 54.245 39.055 ;
    RECT 56.07 38.985 56.34 39.055 ;
    RECT 79.575 38.985 79.645 39.055 ;
    RECT 30.67 38.225 30.74 38.295 ;
    RECT 50.93 38.225 51.0 38.295 ;
    RECT 53.975 38.225 54.245 38.295 ;
    RECT 56.07 38.225 56.34 38.295 ;
    RECT 79.575 38.225 79.645 38.295 ;
    RECT 30.67 37.465 30.74 37.535 ;
    RECT 50.93 37.465 51.0 37.535 ;
    RECT 53.975 37.465 54.245 37.535 ;
    RECT 56.07 37.465 56.34 37.535 ;
    RECT 79.575 37.465 79.645 37.535 ;
    RECT 30.67 36.705 30.74 36.775 ;
    RECT 50.93 36.705 51.0 36.775 ;
    RECT 53.975 36.705 54.245 36.775 ;
    RECT 56.07 36.705 56.34 36.775 ;
    RECT 79.575 36.705 79.645 36.775 ;
    RECT 30.67 35.945 30.74 36.015 ;
    RECT 50.93 35.945 51.0 36.015 ;
    RECT 53.975 35.945 54.245 36.015 ;
    RECT 56.07 35.945 56.34 36.015 ;
    RECT 79.575 35.945 79.645 36.015 ;
    RECT 30.67 35.185 30.74 35.255 ;
    RECT 50.93 35.185 51.0 35.255 ;
    RECT 53.975 35.185 54.245 35.255 ;
    RECT 56.07 35.185 56.34 35.255 ;
    RECT 79.575 35.185 79.645 35.255 ;
    RECT 30.67 34.425 30.74 34.495 ;
    RECT 50.93 34.425 51.0 34.495 ;
    RECT 53.975 34.425 54.245 34.495 ;
    RECT 56.07 34.425 56.34 34.495 ;
    RECT 79.575 34.425 79.645 34.495 ;
    RECT 30.67 33.665 30.74 33.735 ;
    RECT 50.93 33.665 51.0 33.735 ;
    RECT 53.975 33.665 54.245 33.735 ;
    RECT 56.07 33.665 56.34 33.735 ;
    RECT 79.575 33.665 79.645 33.735 ;
    RECT 30.67 32.905 30.74 32.975 ;
    RECT 50.93 32.905 51.0 32.975 ;
    RECT 53.975 32.905 54.245 32.975 ;
    RECT 56.07 32.905 56.34 32.975 ;
    RECT 79.575 32.905 79.645 32.975 ;
    RECT 30.67 32.145 30.74 32.215 ;
    RECT 50.93 32.145 51.0 32.215 ;
    RECT 53.975 32.145 54.245 32.215 ;
    RECT 56.07 32.145 56.34 32.215 ;
    RECT 79.575 32.145 79.645 32.215 ;
    RECT 30.67 31.385 30.74 31.455 ;
    RECT 50.93 31.385 51.0 31.455 ;
    RECT 53.975 31.385 54.245 31.455 ;
    RECT 56.07 31.385 56.34 31.455 ;
    RECT 79.575 31.385 79.645 31.455 ;
    RECT 30.67 30.625 30.74 30.695 ;
    RECT 50.93 30.625 51.0 30.695 ;
    RECT 53.975 30.625 54.245 30.695 ;
    RECT 56.07 30.625 56.34 30.695 ;
    RECT 79.575 30.625 79.645 30.695 ;
    RECT 30.67 29.865 30.74 29.935 ;
    RECT 50.93 29.865 51.0 29.935 ;
    RECT 53.975 29.865 54.245 29.935 ;
    RECT 56.07 29.865 56.34 29.935 ;
    RECT 79.575 29.865 79.645 29.935 ;
    RECT 30.67 29.105 30.74 29.175 ;
    RECT 50.93 29.105 51.0 29.175 ;
    RECT 53.975 29.105 54.245 29.175 ;
    RECT 56.07 29.105 56.34 29.175 ;
    RECT 79.575 29.105 79.645 29.175 ;
    RECT 30.67 28.345 30.74 28.415 ;
    RECT 50.93 28.345 51.0 28.415 ;
    RECT 53.975 28.345 54.245 28.415 ;
    RECT 56.07 28.345 56.34 28.415 ;
    RECT 79.575 28.345 79.645 28.415 ;
    RECT 30.67 27.585 30.74 27.655 ;
    RECT 50.93 27.585 51.0 27.655 ;
    RECT 53.975 27.585 54.245 27.655 ;
    RECT 56.07 27.585 56.34 27.655 ;
    RECT 79.575 27.585 79.645 27.655 ;
    RECT 30.67 26.825 30.74 26.895 ;
    RECT 50.93 26.825 51.0 26.895 ;
    RECT 53.975 26.825 54.245 26.895 ;
    RECT 56.07 26.825 56.34 26.895 ;
    RECT 79.575 26.825 79.645 26.895 ;
    RECT 30.67 26.065 30.74 26.135 ;
    RECT 50.93 26.065 51.0 26.135 ;
    RECT 53.975 26.065 54.245 26.135 ;
    RECT 56.07 26.065 56.34 26.135 ;
    RECT 79.575 26.065 79.645 26.135 ;
    RECT 30.67 25.305 30.74 25.375 ;
    RECT 50.93 25.305 51.0 25.375 ;
    RECT 53.975 25.305 54.245 25.375 ;
    RECT 56.07 25.305 56.34 25.375 ;
    RECT 79.575 25.305 79.645 25.375 ;
    RECT 30.67 24.545 30.74 24.615 ;
    RECT 50.93 24.545 51.0 24.615 ;
    RECT 53.975 24.545 54.245 24.615 ;
    RECT 56.07 24.545 56.34 24.615 ;
    RECT 79.575 24.545 79.645 24.615 ;
    RECT 30.67 23.785 30.74 23.855 ;
    RECT 50.93 23.785 51.0 23.855 ;
    RECT 53.975 23.785 54.245 23.855 ;
    RECT 56.07 23.785 56.34 23.855 ;
    RECT 79.575 23.785 79.645 23.855 ;
    RECT 82.65 11.005 82.86 11.075 ;
    RECT 81.25 11.005 81.46 11.075 ;
    RECT 63.085 110.815 63.295 111.025 ;
    RECT 57.5 110.815 57.71 111.025 ;
    RECT 1.035 110.86 1.245 110.93 ;
    RECT 19.635 110.86 19.845 110.93 ;
    RECT 22.735 110.86 22.945 110.93 ;
    RECT 13.435 110.86 13.645 110.93 ;
    RECT 16.535 110.86 16.745 110.93 ;
    RECT 4.135 110.86 4.345 110.93 ;
    RECT 7.235 110.86 7.445 110.93 ;
    RECT 10.335 110.86 10.545 110.93 ;
    RECT 20.295 60.132 20.505 60.202 ;
    RECT 21.64 60.385 21.85 60.455 ;
    RECT 20.295 109.758 20.505 109.828 ;
    RECT 20.295 10.752 20.505 10.822 ;
    RECT 21.64 109.505 21.85 109.575 ;
    RECT 21.64 11.005 21.85 11.075 ;
    RECT 20.295 110.315 20.505 110.525 ;
    RECT 20.295 10.055 20.505 10.265 ;
    RECT 7.895 60.132 8.105 60.202 ;
    RECT 9.24 60.385 9.45 60.455 ;
    RECT 7.895 109.758 8.105 109.828 ;
    RECT 7.895 10.752 8.105 10.822 ;
    RECT 9.24 109.505 9.45 109.575 ;
    RECT 9.24 11.005 9.45 11.075 ;
    RECT 7.895 110.315 8.105 110.525 ;
    RECT 7.895 10.055 8.105 10.265 ;
    RECT 10.995 60.132 11.205 60.202 ;
    RECT 12.34 60.385 12.55 60.455 ;
    RECT 10.995 109.758 11.205 109.828 ;
    RECT 10.995 10.752 11.205 10.822 ;
    RECT 12.34 109.505 12.55 109.575 ;
    RECT 12.34 11.005 12.55 11.075 ;
    RECT 10.995 110.315 11.205 110.525 ;
    RECT 10.995 10.055 11.205 10.265 ;
    RECT 14.095 60.132 14.305 60.202 ;
    RECT 15.44 60.385 15.65 60.455 ;
    RECT 14.095 109.758 14.305 109.828 ;
    RECT 14.095 10.752 14.305 10.822 ;
    RECT 15.44 109.505 15.65 109.575 ;
    RECT 15.44 11.005 15.65 11.075 ;
    RECT 14.095 110.315 14.305 110.525 ;
    RECT 14.095 10.055 14.305 10.265 ;
    RECT 17.195 60.132 17.405 60.202 ;
    RECT 18.54 60.385 18.75 60.455 ;
    RECT 17.195 109.758 17.405 109.828 ;
    RECT 17.195 10.752 17.405 10.822 ;
    RECT 18.54 109.505 18.75 109.575 ;
    RECT 18.54 11.005 18.75 11.075 ;
    RECT 17.195 110.315 17.405 110.525 ;
    RECT 17.195 10.055 17.405 10.265 ;
    RECT 4.795 60.132 5.005 60.202 ;
    RECT 6.14 60.385 6.35 60.455 ;
    RECT 4.795 109.758 5.005 109.828 ;
    RECT 4.795 10.752 5.005 10.822 ;
    RECT 6.14 109.505 6.35 109.575 ;
    RECT 6.14 11.005 6.35 11.075 ;
    RECT 4.795 110.315 5.005 110.525 ;
    RECT 4.795 10.055 5.005 10.265 ;
    RECT 23.395 60.132 23.605 60.202 ;
    RECT 24.74 60.385 24.95 60.455 ;
    RECT 23.395 109.758 23.605 109.828 ;
    RECT 23.395 10.752 23.605 10.822 ;
    RECT 24.74 109.505 24.95 109.575 ;
    RECT 24.74 11.005 24.95 11.075 ;
    RECT 23.395 110.315 23.605 110.525 ;
    RECT 23.395 10.055 23.605 10.265 ;
    RECT 1.695 60.132 1.905 60.202 ;
    RECT 3.04 60.385 3.25 60.455 ;
    RECT 1.695 109.758 1.905 109.828 ;
    RECT 1.695 10.752 1.905 10.822 ;
    RECT 3.04 109.505 3.25 109.575 ;
    RECT 3.04 11.005 3.25 11.075 ;
    RECT 1.695 110.315 1.905 110.525 ;
    RECT 1.695 10.055 1.905 10.265 ;
    RECT 0.77 3.27 0.84 3.34 ;
    RECT 0.76 2.545 0.83 2.615 ;
    RECT 0.755 9.475 0.825 9.685 ;
    RECT 0.77 8.1 0.84 8.17 ;
    RECT 13.435 0.645 13.645 0.715 ;
    RECT 16.535 0.645 16.745 0.715 ;
    RECT 19.635 0.645 19.845 0.715 ;
    RECT 22.735 0.645 22.945 0.715 ;
    RECT 1.035 0.645 1.245 0.715 ;
    RECT 4.135 0.645 4.345 0.715 ;
    RECT 7.235 0.645 7.445 0.715 ;
    RECT 10.335 0.645 10.545 0.715 ;
    RECT 6.14 1.375 6.35 1.585 ;
    RECT 9.895 2.01 10.105 2.08 ;
    RECT 12.995 2.01 13.205 2.08 ;
    RECT 15.44 1.375 15.65 1.585 ;
    RECT 16.535 2.52 16.745 2.59 ;
    RECT 18.54 1.375 18.75 1.585 ;
    RECT 22.295 2.01 22.505 2.08 ;
    RECT 25.395 2.01 25.605 2.08 ;
    RECT 9.24 1.375 9.45 1.585 ;
    RECT 10.335 2.52 10.545 2.59 ;
    RECT 3.695 2.01 3.905 2.08 ;
    RECT 6.795 2.01 7.005 2.08 ;
    RECT 12.34 1.375 12.55 1.585 ;
    RECT 16.095 2.01 16.305 2.08 ;
    RECT 21.64 1.375 21.85 1.585 ;
    RECT 22.735 2.52 22.945 2.59 ;
    RECT 24.74 1.375 24.95 1.585 ;
    RECT 19.195 2.01 19.405 2.08 ;
    RECT 3.04 1.375 3.25 1.585 ;
    RECT 4.135 2.52 4.345 2.59 ;
    RECT 21.64 7.09 21.85 7.16 ;
    RECT 21.64 3.65 21.85 3.72 ;
    RECT 21.64 2.86 21.85 2.93 ;
    RECT 24.74 7.09 24.95 7.16 ;
    RECT 24.74 3.65 24.95 3.72 ;
    RECT 24.74 2.86 24.95 2.93 ;
    RECT 3.04 6.31 3.25 6.38 ;
    RECT 6.14 6.31 6.35 6.38 ;
    RECT 3.695 4.72 3.905 4.79 ;
    RECT 6.795 4.72 7.005 4.79 ;
    RECT 3.04 7.09 3.25 7.16 ;
    RECT 3.04 3.65 3.25 3.72 ;
    RECT 3.04 2.86 3.25 2.93 ;
    RECT 12.995 4.72 13.205 4.79 ;
    RECT 9.24 7.09 9.45 7.16 ;
    RECT 9.24 3.65 9.45 3.72 ;
    RECT 9.24 2.86 9.45 2.93 ;
    RECT 6.14 7.09 6.35 7.16 ;
    RECT 12.34 7.09 12.55 7.16 ;
    RECT 6.14 3.65 6.35 3.72 ;
    RECT 12.34 3.65 12.55 3.72 ;
    RECT 6.14 2.86 6.35 2.93 ;
    RECT 12.34 2.86 12.55 2.93 ;
    RECT 15.44 6.31 15.65 6.38 ;
    RECT 9.24 6.31 9.45 6.38 ;
    RECT 12.34 6.31 12.55 6.38 ;
    RECT 9.895 4.72 10.105 4.79 ;
    RECT 18.54 6.31 18.75 6.38 ;
    RECT 16.095 4.72 16.305 4.79 ;
    RECT 19.195 4.72 19.405 4.79 ;
    RECT 15.44 7.09 15.65 7.16 ;
    RECT 15.44 3.65 15.65 3.72 ;
    RECT 15.44 2.86 15.65 2.93 ;
    RECT 18.54 7.09 18.75 7.16 ;
    RECT 18.54 3.65 18.75 3.72 ;
    RECT 18.54 2.86 18.75 2.93 ;
    RECT 21.64 6.31 21.85 6.38 ;
    RECT 24.74 6.31 24.95 6.38 ;
    RECT 22.295 4.72 22.505 4.79 ;
    RECT 25.395 4.72 25.605 4.79 ;
    RECT 96.57 0.645 96.78 0.715 ;
    RECT 93.47 0.645 93.68 0.715 ;
    RECT 90.37 0.645 90.58 0.715 ;
    RECT 87.27 0.645 87.48 0.715 ;
    RECT 108.97 0.645 109.18 0.715 ;
    RECT 105.87 0.645 106.08 0.715 ;
    RECT 102.77 0.645 102.98 0.715 ;
    RECT 99.67 0.645 99.88 0.715 ;
    RECT 84.61 2.01 84.82 2.08 ;
    RECT 97.665 1.375 97.875 1.585 ;
    RECT 88.365 1.375 88.575 1.585 ;
    RECT 87.27 2.52 87.48 2.59 ;
    RECT 85.265 1.375 85.475 1.585 ;
    RECT 106.965 1.375 107.175 1.585 ;
    RECT 105.87 2.52 106.08 2.59 ;
    RECT 103.865 1.375 104.075 1.585 ;
    RECT 106.31 2.01 106.52 2.08 ;
    RECT 103.21 2.01 103.42 2.08 ;
    RECT 93.91 2.01 94.12 2.08 ;
    RECT 90.81 2.01 91.02 2.08 ;
    RECT 94.565 1.375 94.775 1.585 ;
    RECT 93.47 2.52 93.68 2.59 ;
    RECT 91.465 1.375 91.675 1.585 ;
    RECT 100.11 2.01 100.32 2.08 ;
    RECT 97.01 2.01 97.22 2.08 ;
    RECT 87.71 2.01 87.92 2.08 ;
    RECT 100.765 1.375 100.975 1.585 ;
    RECT 99.67 2.52 99.88 2.59 ;
    RECT 88.365 7.09 88.575 7.16 ;
    RECT 88.365 3.65 88.575 3.72 ;
    RECT 106.965 6.31 107.175 6.38 ;
    RECT 103.865 6.31 104.075 6.38 ;
    RECT 88.365 2.86 88.575 2.93 ;
    RECT 85.265 7.09 85.475 7.16 ;
    RECT 85.265 3.65 85.475 3.72 ;
    RECT 85.265 2.86 85.475 2.93 ;
    RECT 106.31 4.72 106.52 4.79 ;
    RECT 103.21 4.72 103.42 4.79 ;
    RECT 106.965 7.09 107.175 7.16 ;
    RECT 106.965 3.65 107.175 3.72 ;
    RECT 106.965 2.86 107.175 2.93 ;
    RECT 103.865 7.09 104.075 7.16 ;
    RECT 103.865 3.65 104.075 3.72 ;
    RECT 103.865 2.86 104.075 2.93 ;
    RECT 100.765 6.31 100.975 6.38 ;
    RECT 97.665 6.31 97.875 6.38 ;
    RECT 100.11 4.72 100.32 4.79 ;
    RECT 97.01 4.72 97.22 4.79 ;
    RECT 100.765 7.09 100.975 7.16 ;
    RECT 100.765 3.65 100.975 3.72 ;
    RECT 100.765 2.86 100.975 2.93 ;
    RECT 97.665 7.09 97.875 7.16 ;
    RECT 97.665 3.65 97.875 3.72 ;
    RECT 97.665 2.86 97.875 2.93 ;
    RECT 94.565 6.31 94.775 6.38 ;
    RECT 91.465 6.31 91.675 6.38 ;
    RECT 93.91 4.72 94.12 4.79 ;
    RECT 90.81 4.72 91.02 4.79 ;
    RECT 94.565 7.09 94.775 7.16 ;
    RECT 94.565 3.65 94.775 3.72 ;
    RECT 94.565 2.86 94.775 2.93 ;
    RECT 91.465 7.09 91.675 7.16 ;
    RECT 91.465 3.65 91.675 3.72 ;
    RECT 91.465 2.86 91.675 2.93 ;
    RECT 88.365 6.31 88.575 6.38 ;
    RECT 85.265 6.31 85.475 6.38 ;
    RECT 87.71 4.72 87.92 4.79 ;
    RECT 84.61 4.72 84.82 4.79 ;
    RECT 109.39 9.475 109.46 9.685 ;
    RECT 109.385 2.545 109.455 2.615 ;
    RECT 109.375 8.1 109.445 8.17 ;
    RECT 109.375 3.27 109.445 3.34 ;
    LAYER M4 DESIGNRULEWIDTH 0.165 ;
    RECT 26.78 0.0 27.32 0.78 ;
    RECT 27.8 0.0 28.02 0.78 ;
    RECT 28.5 0.0 28.72 0.78 ;
    RECT 29.2 0.0 30.815 0.78 ;
    RECT 31.295 0.0 31.515 0.78 ;
    RECT 31.995 0.0 32.21 0.78 ;
    RECT 32.69 0.0 32.91 0.78 ;
    RECT 33.39 0.0 33.61 0.78 ;
    RECT 34.09 0.0 34.31 0.78 ;
    RECT 34.79 0.0 35.005 0.78 ;
    RECT 35.485 0.32 36.405 0.78 ;
    RECT 35.485 0.0 35.75 0.32 ;
    RECT 36.17 0.0 36.405 0.32 ;
    RECT 36.885 0.0 37.105 0.78 ;
    RECT 37.585 0.0 37.8 0.78 ;
    RECT 38.28 0.0 38.5 0.78 ;
    RECT 38.98 0.0 39.2 0.78 ;
    RECT 39.68 0.0 39.895 0.78 ;
    RECT 40.375 0.0 40.595 0.78 ;
    RECT 41.075 0.0 41.995 0.78 ;
    RECT 42.475 0.0 42.69 0.78 ;
    RECT 43.17 0.0 43.39 0.78 ;
    RECT 43.87 0.0 44.09 0.78 ;
    RECT 44.57 0.0 44.79 0.78 ;
    RECT 45.27 0.32 45.485 0.78 ;
    RECT 45.965 0.0 46.185 0.78 ;
    RECT 46.665 0.0 47.58 0.78 ;
    RECT 48.06 0.0 48.28 0.78 ;
    RECT 48.76 0.0 48.98 0.78 ;
    RECT 49.46 0.0 49.68 0.78 ;
    RECT 50.16 0.0 50.375 0.78 ;
    RECT 50.855 0.0 51.775 0.78 ;
    RECT 52.255 0.0 53.17 0.78 ;
    RECT 53.65 0.0 53.87 0.78 ;
    RECT 54.35 0.0 54.57 0.78 ;
    RECT 55.05 0.0 55.265 0.78 ;
    RECT 55.745 0.0 55.965 0.78 ;
    RECT 56.445 0.0 56.665 0.78 ;
    RECT 57.145 0.0 58.06 0.78 ;
    RECT 58.54 0.0 59.46 0.78 ;
    RECT 59.94 0.0 60.16 0.78 ;
    RECT 60.64 0.0 60.855 0.78 ;
    RECT 61.335 0.0 61.555 0.78 ;
    RECT 62.035 0.0 62.25 0.78 ;
    RECT 62.73 0.0 63.65 0.78 ;
    RECT 64.13 0.0 64.345 0.78 ;
    RECT 64.825 0.0 65.045 0.78 ;
    RECT 65.525 0.0 65.745 0.78 ;
    RECT 66.225 0.0 66.445 0.78 ;
    RECT 66.925 0.0 67.14 0.78 ;
    RECT 67.62 0.0 67.84 0.78 ;
    RECT 68.32 0.0 69.235 0.78 ;
    RECT 69.715 0.0 69.935 0.78 ;
    RECT 70.415 0.0 70.635 0.78 ;
    RECT 71.115 0.0 71.335 0.78 ;
    RECT 71.815 0.0 72.035 0.78 ;
    RECT 72.515 0.0 72.735 0.78 ;
    RECT 73.215 0.0 73.435 0.78 ;
    RECT 73.915 0.0 74.835 0.78 ;
    RECT 75.315 0.0 75.535 0.78 ;
    RECT 76.015 0.0 76.225 0.36 ;
    RECT 76.705 0.0 76.92 0.36 ;
    RECT 77.4 0.0 77.62 0.78 ;
    RECT 78.1 0.0 78.32 0.78 ;
    RECT 78.8 0.0 79.02 0.78 ;
    RECT 79.5 0.0 81.115 0.78 ;
    RECT 81.595 0.0 81.815 0.78 ;
    RECT 82.295 0.0 82.515 0.78 ;
    RECT 82.995 0.0 83.435 0.78 ;
    RECT 26.78 0.78 27.32 9.81 ;
    RECT 27.8 0.78 28.02 9.81 ;
    RECT 28.5 0.78 28.72 9.81 ;
    RECT 29.2 0.78 30.815 9.81 ;
    RECT 31.295 0.78 31.515 9.81 ;
    RECT 31.995 0.78 32.21 9.81 ;
    RECT 32.69 0.78 32.91 9.81 ;
    RECT 33.39 0.78 33.61 9.81 ;
    RECT 34.09 0.78 34.31 9.81 ;
    RECT 34.79 0.78 35.005 9.81 ;
    RECT 35.485 0.78 36.405 9.81 ;
    RECT 36.885 0.78 37.105 9.81 ;
    RECT 37.585 0.78 37.8 9.81 ;
    RECT 38.28 0.78 38.5 9.81 ;
    RECT 38.98 0.78 39.2 9.81 ;
    RECT 39.68 0.78 39.895 9.81 ;
    RECT 40.375 0.78 40.595 9.81 ;
    RECT 41.075 0.78 41.995 9.81 ;
    RECT 42.475 0.78 42.69 9.81 ;
    RECT 43.17 0.78 43.39 9.81 ;
    RECT 43.87 0.78 44.09 9.81 ;
    RECT 44.57 0.78 44.79 9.81 ;
    RECT 45.27 0.78 45.485 9.81 ;
    RECT 45.965 0.78 46.185 9.81 ;
    RECT 46.665 0.78 47.58 9.81 ;
    RECT 48.06 0.78 48.28 9.81 ;
    RECT 48.76 0.78 48.98 9.81 ;
    RECT 49.46 0.78 49.68 9.81 ;
    RECT 50.16 0.78 50.375 9.81 ;
    RECT 50.855 0.78 51.775 9.81 ;
    RECT 52.255 0.78 53.17 9.81 ;
    RECT 53.65 0.78 53.87 1.795 ;
    RECT 53.65 9.555 53.87 9.81 ;
    RECT 54.35 0.78 54.57 9.81 ;
    RECT 55.05 0.78 55.265 9.81 ;
    RECT 55.745 0.78 55.965 9.81 ;
    RECT 56.445 0.78 56.665 9.81 ;
    RECT 57.145 0.78 58.06 9.81 ;
    RECT 58.54 0.78 59.46 9.81 ;
    RECT 59.94 0.78 60.16 9.81 ;
    RECT 60.64 0.78 60.855 9.81 ;
    RECT 61.335 0.78 61.555 9.81 ;
    RECT 62.035 0.78 62.25 9.81 ;
    RECT 62.73 0.78 63.65 9.81 ;
    RECT 64.13 0.78 64.345 9.81 ;
    RECT 64.825 0.78 65.045 9.81 ;
    RECT 65.525 0.78 65.745 9.81 ;
    RECT 66.225 0.78 66.445 9.81 ;
    RECT 66.925 0.78 67.14 9.81 ;
    RECT 67.62 0.78 67.84 9.81 ;
    RECT 68.32 0.78 69.235 9.81 ;
    RECT 69.715 0.78 69.935 9.81 ;
    RECT 70.415 0.78 70.635 9.81 ;
    RECT 71.115 0.78 71.335 9.81 ;
    RECT 71.815 0.78 72.035 9.81 ;
    RECT 72.515 0.78 72.735 9.81 ;
    RECT 73.215 0.78 73.435 9.81 ;
    RECT 73.915 0.78 74.6 9.81 ;
    RECT 74.6 1.305 74.835 9.81 ;
    RECT 75.315 0.78 75.535 9.81 ;
    RECT 76.015 0.78 76.225 9.81 ;
    RECT 76.705 0.78 76.92 9.81 ;
    RECT 77.4 0.78 77.62 9.81 ;
    RECT 78.1 0.78 78.32 9.81 ;
    RECT 78.8 0.78 79.02 9.81 ;
    RECT 79.5 0.78 81.115 9.81 ;
    RECT 81.595 0.78 81.815 9.81 ;
    RECT 82.295 0.78 82.515 9.81 ;
    RECT 82.995 0.78 83.435 9.81 ;
    RECT 105.835 110.77 106.115 110.975 ;
    RECT 102.735 110.77 103.015 110.975 ;
    RECT 99.635 110.77 99.915 110.975 ;
    RECT 96.535 110.77 96.815 110.975 ;
    RECT 93.435 110.77 93.715 110.975 ;
    RECT 90.335 110.77 90.615 110.975 ;
    RECT 87.235 110.77 87.515 110.975 ;
    RECT 108.935 110.77 109.215 110.975 ;
    RECT 90.335 31.8 90.615 32.56 ;
    RECT 90.335 31.04 90.615 31.8 ;
    RECT 90.335 30.28 90.615 31.04 ;
    RECT 90.335 29.52 90.615 30.28 ;
    RECT 90.335 28.76 90.615 29.52 ;
    RECT 90.335 28.0 90.615 28.76 ;
    RECT 90.335 27.24 90.615 28.0 ;
    RECT 90.335 26.48 90.615 27.24 ;
    RECT 90.335 100.18 90.615 100.94 ;
    RECT 90.335 25.72 90.615 26.48 ;
    RECT 90.335 99.42 90.615 100.18 ;
    RECT 90.335 24.96 90.615 25.72 ;
    RECT 90.335 98.66 90.615 99.42 ;
    RECT 90.335 97.9 90.615 98.66 ;
    RECT 90.335 97.14 90.615 97.9 ;
    RECT 90.335 96.38 90.615 97.14 ;
    RECT 90.335 95.62 90.615 96.38 ;
    RECT 90.335 94.86 90.615 95.62 ;
    RECT 90.335 94.1 90.615 94.86 ;
    RECT 90.335 93.34 90.615 94.1 ;
    RECT 90.335 24.2 90.615 24.96 ;
    RECT 90.335 23.44 90.615 24.2 ;
    RECT 90.335 22.68 90.615 23.44 ;
    RECT 90.335 21.92 90.615 22.68 ;
    RECT 90.335 21.16 90.615 21.92 ;
    RECT 90.335 20.4 90.615 21.16 ;
    RECT 90.335 19.64 90.615 20.4 ;
    RECT 90.335 18.88 90.615 19.64 ;
    RECT 90.335 92.58 90.615 93.34 ;
    RECT 90.335 18.12 90.615 18.88 ;
    RECT 90.335 91.82 90.615 92.58 ;
    RECT 90.335 17.36 90.615 18.12 ;
    RECT 90.335 91.06 90.615 91.82 ;
    RECT 90.335 90.3 90.615 91.06 ;
    RECT 90.335 89.54 90.615 90.3 ;
    RECT 90.335 88.78 90.615 89.54 ;
    RECT 90.335 88.02 90.615 88.78 ;
    RECT 90.335 87.26 90.615 88.02 ;
    RECT 90.335 86.5 90.615 87.26 ;
    RECT 90.335 85.74 90.615 86.5 ;
    RECT 90.335 84.98 90.615 85.74 ;
    RECT 90.335 84.22 90.615 84.98 ;
    RECT 90.335 83.46 90.615 84.22 ;
    RECT 90.335 82.7 90.615 83.46 ;
    RECT 90.335 81.94 90.615 82.7 ;
    RECT 90.335 81.18 90.615 81.94 ;
    RECT 90.335 80.42 90.615 81.18 ;
    RECT 90.335 79.66 90.615 80.42 ;
    RECT 90.335 78.9 90.615 79.66 ;
    RECT 90.335 78.14 90.615 78.9 ;
    RECT 90.335 77.38 90.615 78.14 ;
    RECT 90.335 76.62 90.615 77.38 ;
    RECT 90.335 75.86 90.615 76.62 ;
    RECT 90.335 75.1 90.615 75.86 ;
    RECT 90.335 74.34 90.615 75.1 ;
    RECT 90.335 73.58 90.615 74.34 ;
    RECT 90.335 72.82 90.615 73.58 ;
    RECT 90.335 72.06 90.615 72.82 ;
    RECT 90.335 71.3 90.615 72.06 ;
    RECT 90.335 70.54 90.615 71.3 ;
    RECT 90.335 69.78 90.615 70.54 ;
    RECT 90.335 69.02 90.615 69.78 ;
    RECT 90.335 68.26 90.615 69.02 ;
    RECT 90.335 67.5 90.615 68.26 ;
    RECT 90.335 66.74 90.615 67.5 ;
    RECT 90.335 65.98 90.615 66.74 ;
    RECT 90.335 65.22 90.615 65.98 ;
    RECT 90.335 64.46 90.615 65.22 ;
    RECT 90.335 63.7 90.615 64.46 ;
    RECT 90.335 62.94 90.615 63.7 ;
    RECT 90.335 108.54 90.615 109.3 ;
    RECT 90.335 62.18 90.615 62.94 ;
    RECT 90.335 61.42 90.615 62.18 ;
    RECT 90.335 60.66 90.615 61.42 ;
    RECT 90.335 59.92 90.615 60.66 ;
    RECT 90.335 59.16 90.615 59.92 ;
    RECT 90.335 58.4 90.615 59.16 ;
    RECT 90.335 57.64 90.615 58.4 ;
    RECT 90.335 56.88 90.615 57.64 ;
    RECT 90.335 56.12 90.615 56.88 ;
    RECT 90.335 55.36 90.615 56.12 ;
    RECT 90.335 16.6 90.615 17.36 ;
    RECT 90.335 15.84 90.615 16.6 ;
    RECT 90.335 15.08 90.615 15.84 ;
    RECT 90.335 14.32 90.615 15.08 ;
    RECT 90.335 13.56 90.615 14.32 ;
    RECT 90.335 12.8 90.615 13.56 ;
    RECT 90.335 12.04 90.615 12.8 ;
    RECT 90.335 9.81 90.615 11.28 ;
    RECT 90.335 54.6 90.615 55.36 ;
    RECT 90.335 53.84 90.615 54.6 ;
    RECT 90.335 53.08 90.615 53.84 ;
    RECT 90.335 52.32 90.615 53.08 ;
    RECT 90.335 51.56 90.615 52.32 ;
    RECT 90.335 50.8 90.615 51.56 ;
    RECT 90.335 50.04 90.615 50.8 ;
    RECT 90.335 49.28 90.615 50.04 ;
    RECT 90.335 48.52 90.615 49.28 ;
    RECT 90.335 47.76 90.615 48.52 ;
    RECT 90.335 11.28 90.615 12.04 ;
    RECT 90.335 47.0 90.615 47.76 ;
    RECT 90.335 46.24 90.615 47.0 ;
    RECT 90.335 45.48 90.615 46.24 ;
    RECT 90.335 44.72 90.615 45.48 ;
    RECT 90.335 43.96 90.615 44.72 ;
    RECT 90.335 43.2 90.615 43.96 ;
    RECT 90.335 42.44 90.615 43.2 ;
    RECT 90.335 41.68 90.615 42.44 ;
    RECT 90.335 40.92 90.615 41.68 ;
    RECT 90.335 40.16 90.615 40.92 ;
    RECT 90.335 109.3 90.615 110.77 ;
    RECT 90.335 39.4 90.615 40.16 ;
    RECT 90.335 38.64 90.615 39.4 ;
    RECT 90.335 37.88 90.615 38.64 ;
    RECT 90.335 37.12 90.615 37.88 ;
    RECT 90.335 36.36 90.615 37.12 ;
    RECT 90.335 35.6 90.615 36.36 ;
    RECT 90.335 34.84 90.615 35.6 ;
    RECT 90.335 34.08 90.615 34.84 ;
    RECT 90.335 107.78 90.615 108.54 ;
    RECT 90.335 33.32 90.615 34.08 ;
    RECT 90.335 107.02 90.615 107.78 ;
    RECT 90.335 32.56 90.615 33.32 ;
    RECT 90.335 106.26 90.615 107.02 ;
    RECT 90.335 105.5 90.615 106.26 ;
    RECT 90.335 104.74 90.615 105.5 ;
    RECT 90.335 103.98 90.615 104.74 ;
    RECT 90.335 103.22 90.615 103.98 ;
    RECT 90.335 102.46 90.615 103.22 ;
    RECT 90.335 101.7 90.615 102.46 ;
    RECT 90.335 100.94 90.615 101.7 ;
    RECT 102.735 31.8 103.015 32.56 ;
    RECT 102.735 31.04 103.015 31.8 ;
    RECT 102.735 30.28 103.015 31.04 ;
    RECT 102.735 29.52 103.015 30.28 ;
    RECT 102.735 28.76 103.015 29.52 ;
    RECT 102.735 28.0 103.015 28.76 ;
    RECT 102.735 27.24 103.015 28.0 ;
    RECT 102.735 26.48 103.015 27.24 ;
    RECT 102.735 100.18 103.015 100.94 ;
    RECT 102.735 25.72 103.015 26.48 ;
    RECT 102.735 99.42 103.015 100.18 ;
    RECT 102.735 24.96 103.015 25.72 ;
    RECT 102.735 98.66 103.015 99.42 ;
    RECT 102.735 97.9 103.015 98.66 ;
    RECT 102.735 97.14 103.015 97.9 ;
    RECT 102.735 96.38 103.015 97.14 ;
    RECT 102.735 95.62 103.015 96.38 ;
    RECT 102.735 94.86 103.015 95.62 ;
    RECT 102.735 94.1 103.015 94.86 ;
    RECT 102.735 93.34 103.015 94.1 ;
    RECT 102.735 24.2 103.015 24.96 ;
    RECT 102.735 23.44 103.015 24.2 ;
    RECT 102.735 22.68 103.015 23.44 ;
    RECT 102.735 21.92 103.015 22.68 ;
    RECT 102.735 21.16 103.015 21.92 ;
    RECT 102.735 20.4 103.015 21.16 ;
    RECT 102.735 19.64 103.015 20.4 ;
    RECT 102.735 18.88 103.015 19.64 ;
    RECT 102.735 92.58 103.015 93.34 ;
    RECT 102.735 18.12 103.015 18.88 ;
    RECT 102.735 91.82 103.015 92.58 ;
    RECT 102.735 17.36 103.015 18.12 ;
    RECT 102.735 91.06 103.015 91.82 ;
    RECT 102.735 90.3 103.015 91.06 ;
    RECT 102.735 89.54 103.015 90.3 ;
    RECT 102.735 88.78 103.015 89.54 ;
    RECT 102.735 88.02 103.015 88.78 ;
    RECT 102.735 87.26 103.015 88.02 ;
    RECT 102.735 86.5 103.015 87.26 ;
    RECT 102.735 85.74 103.015 86.5 ;
    RECT 102.735 84.98 103.015 85.74 ;
    RECT 102.735 84.22 103.015 84.98 ;
    RECT 102.735 83.46 103.015 84.22 ;
    RECT 102.735 82.7 103.015 83.46 ;
    RECT 102.735 81.94 103.015 82.7 ;
    RECT 102.735 81.18 103.015 81.94 ;
    RECT 102.735 80.42 103.015 81.18 ;
    RECT 102.735 79.66 103.015 80.42 ;
    RECT 102.735 78.9 103.015 79.66 ;
    RECT 102.735 78.14 103.015 78.9 ;
    RECT 102.735 77.38 103.015 78.14 ;
    RECT 102.735 76.62 103.015 77.38 ;
    RECT 102.735 75.86 103.015 76.62 ;
    RECT 102.735 75.1 103.015 75.86 ;
    RECT 102.735 74.34 103.015 75.1 ;
    RECT 102.735 73.58 103.015 74.34 ;
    RECT 102.735 72.82 103.015 73.58 ;
    RECT 102.735 72.06 103.015 72.82 ;
    RECT 102.735 71.3 103.015 72.06 ;
    RECT 102.735 70.54 103.015 71.3 ;
    RECT 102.735 69.78 103.015 70.54 ;
    RECT 102.735 69.02 103.015 69.78 ;
    RECT 102.735 68.26 103.015 69.02 ;
    RECT 102.735 67.5 103.015 68.26 ;
    RECT 102.735 66.74 103.015 67.5 ;
    RECT 102.735 65.98 103.015 66.74 ;
    RECT 102.735 65.22 103.015 65.98 ;
    RECT 102.735 64.46 103.015 65.22 ;
    RECT 102.735 63.7 103.015 64.46 ;
    RECT 102.735 62.94 103.015 63.7 ;
    RECT 102.735 108.54 103.015 109.3 ;
    RECT 102.735 62.18 103.015 62.94 ;
    RECT 102.735 61.42 103.015 62.18 ;
    RECT 102.735 60.66 103.015 61.42 ;
    RECT 102.735 59.92 103.015 60.66 ;
    RECT 102.735 59.16 103.015 59.92 ;
    RECT 102.735 58.4 103.015 59.16 ;
    RECT 102.735 57.64 103.015 58.4 ;
    RECT 102.735 56.88 103.015 57.64 ;
    RECT 102.735 56.12 103.015 56.88 ;
    RECT 102.735 55.36 103.015 56.12 ;
    RECT 102.735 16.6 103.015 17.36 ;
    RECT 102.735 15.84 103.015 16.6 ;
    RECT 102.735 15.08 103.015 15.84 ;
    RECT 102.735 14.32 103.015 15.08 ;
    RECT 102.735 13.56 103.015 14.32 ;
    RECT 102.735 12.8 103.015 13.56 ;
    RECT 102.735 12.04 103.015 12.8 ;
    RECT 102.735 9.81 103.015 11.28 ;
    RECT 102.735 54.6 103.015 55.36 ;
    RECT 102.735 53.84 103.015 54.6 ;
    RECT 102.735 53.08 103.015 53.84 ;
    RECT 102.735 52.32 103.015 53.08 ;
    RECT 102.735 51.56 103.015 52.32 ;
    RECT 102.735 50.8 103.015 51.56 ;
    RECT 102.735 50.04 103.015 50.8 ;
    RECT 102.735 49.28 103.015 50.04 ;
    RECT 102.735 48.52 103.015 49.28 ;
    RECT 102.735 47.76 103.015 48.52 ;
    RECT 102.735 11.28 103.015 12.04 ;
    RECT 102.735 47.0 103.015 47.76 ;
    RECT 102.735 46.24 103.015 47.0 ;
    RECT 102.735 45.48 103.015 46.24 ;
    RECT 102.735 44.72 103.015 45.48 ;
    RECT 102.735 43.96 103.015 44.72 ;
    RECT 102.735 43.2 103.015 43.96 ;
    RECT 102.735 42.44 103.015 43.2 ;
    RECT 102.735 41.68 103.015 42.44 ;
    RECT 102.735 40.92 103.015 41.68 ;
    RECT 102.735 40.16 103.015 40.92 ;
    RECT 102.735 109.3 103.015 110.77 ;
    RECT 102.735 39.4 103.015 40.16 ;
    RECT 102.735 38.64 103.015 39.4 ;
    RECT 102.735 37.88 103.015 38.64 ;
    RECT 102.735 37.12 103.015 37.88 ;
    RECT 102.735 36.36 103.015 37.12 ;
    RECT 102.735 35.6 103.015 36.36 ;
    RECT 102.735 34.84 103.015 35.6 ;
    RECT 102.735 34.08 103.015 34.84 ;
    RECT 102.735 107.78 103.015 108.54 ;
    RECT 102.735 33.32 103.015 34.08 ;
    RECT 102.735 107.02 103.015 107.78 ;
    RECT 102.735 32.56 103.015 33.32 ;
    RECT 102.735 106.26 103.015 107.02 ;
    RECT 102.735 105.5 103.015 106.26 ;
    RECT 102.735 104.74 103.015 105.5 ;
    RECT 102.735 103.98 103.015 104.74 ;
    RECT 102.735 103.22 103.015 103.98 ;
    RECT 102.735 102.46 103.015 103.22 ;
    RECT 102.735 101.7 103.015 102.46 ;
    RECT 102.735 100.94 103.015 101.7 ;
    RECT 99.635 31.8 99.915 32.56 ;
    RECT 99.635 31.04 99.915 31.8 ;
    RECT 99.635 30.28 99.915 31.04 ;
    RECT 99.635 29.52 99.915 30.28 ;
    RECT 99.635 28.76 99.915 29.52 ;
    RECT 99.635 28.0 99.915 28.76 ;
    RECT 99.635 27.24 99.915 28.0 ;
    RECT 99.635 26.48 99.915 27.24 ;
    RECT 99.635 100.18 99.915 100.94 ;
    RECT 99.635 25.72 99.915 26.48 ;
    RECT 99.635 99.42 99.915 100.18 ;
    RECT 99.635 24.96 99.915 25.72 ;
    RECT 99.635 98.66 99.915 99.42 ;
    RECT 99.635 97.9 99.915 98.66 ;
    RECT 99.635 97.14 99.915 97.9 ;
    RECT 99.635 96.38 99.915 97.14 ;
    RECT 99.635 95.62 99.915 96.38 ;
    RECT 99.635 94.86 99.915 95.62 ;
    RECT 99.635 94.1 99.915 94.86 ;
    RECT 99.635 93.34 99.915 94.1 ;
    RECT 99.635 24.2 99.915 24.96 ;
    RECT 99.635 23.44 99.915 24.2 ;
    RECT 99.635 22.68 99.915 23.44 ;
    RECT 99.635 21.92 99.915 22.68 ;
    RECT 99.635 21.16 99.915 21.92 ;
    RECT 99.635 20.4 99.915 21.16 ;
    RECT 99.635 19.64 99.915 20.4 ;
    RECT 99.635 18.88 99.915 19.64 ;
    RECT 99.635 92.58 99.915 93.34 ;
    RECT 99.635 18.12 99.915 18.88 ;
    RECT 99.635 91.82 99.915 92.58 ;
    RECT 99.635 17.36 99.915 18.12 ;
    RECT 99.635 91.06 99.915 91.82 ;
    RECT 99.635 90.3 99.915 91.06 ;
    RECT 99.635 89.54 99.915 90.3 ;
    RECT 99.635 88.78 99.915 89.54 ;
    RECT 99.635 88.02 99.915 88.78 ;
    RECT 99.635 87.26 99.915 88.02 ;
    RECT 99.635 86.5 99.915 87.26 ;
    RECT 99.635 85.74 99.915 86.5 ;
    RECT 99.635 84.98 99.915 85.74 ;
    RECT 99.635 84.22 99.915 84.98 ;
    RECT 99.635 83.46 99.915 84.22 ;
    RECT 99.635 82.7 99.915 83.46 ;
    RECT 99.635 81.94 99.915 82.7 ;
    RECT 99.635 81.18 99.915 81.94 ;
    RECT 99.635 80.42 99.915 81.18 ;
    RECT 99.635 79.66 99.915 80.42 ;
    RECT 99.635 78.9 99.915 79.66 ;
    RECT 99.635 78.14 99.915 78.9 ;
    RECT 99.635 77.38 99.915 78.14 ;
    RECT 99.635 76.62 99.915 77.38 ;
    RECT 99.635 75.86 99.915 76.62 ;
    RECT 99.635 75.1 99.915 75.86 ;
    RECT 99.635 74.34 99.915 75.1 ;
    RECT 99.635 73.58 99.915 74.34 ;
    RECT 99.635 72.82 99.915 73.58 ;
    RECT 99.635 72.06 99.915 72.82 ;
    RECT 99.635 71.3 99.915 72.06 ;
    RECT 99.635 70.54 99.915 71.3 ;
    RECT 99.635 69.78 99.915 70.54 ;
    RECT 99.635 69.02 99.915 69.78 ;
    RECT 99.635 68.26 99.915 69.02 ;
    RECT 99.635 67.5 99.915 68.26 ;
    RECT 99.635 66.74 99.915 67.5 ;
    RECT 99.635 65.98 99.915 66.74 ;
    RECT 99.635 65.22 99.915 65.98 ;
    RECT 99.635 64.46 99.915 65.22 ;
    RECT 99.635 63.7 99.915 64.46 ;
    RECT 99.635 62.94 99.915 63.7 ;
    RECT 99.635 108.54 99.915 109.3 ;
    RECT 99.635 62.18 99.915 62.94 ;
    RECT 99.635 61.42 99.915 62.18 ;
    RECT 99.635 60.66 99.915 61.42 ;
    RECT 99.635 59.92 99.915 60.66 ;
    RECT 99.635 59.16 99.915 59.92 ;
    RECT 99.635 58.4 99.915 59.16 ;
    RECT 99.635 57.64 99.915 58.4 ;
    RECT 99.635 56.88 99.915 57.64 ;
    RECT 99.635 56.12 99.915 56.88 ;
    RECT 99.635 55.36 99.915 56.12 ;
    RECT 99.635 16.6 99.915 17.36 ;
    RECT 99.635 15.84 99.915 16.6 ;
    RECT 99.635 15.08 99.915 15.84 ;
    RECT 99.635 14.32 99.915 15.08 ;
    RECT 99.635 13.56 99.915 14.32 ;
    RECT 99.635 12.8 99.915 13.56 ;
    RECT 99.635 12.04 99.915 12.8 ;
    RECT 99.635 9.81 99.915 11.28 ;
    RECT 99.635 54.6 99.915 55.36 ;
    RECT 99.635 53.84 99.915 54.6 ;
    RECT 99.635 53.08 99.915 53.84 ;
    RECT 99.635 52.32 99.915 53.08 ;
    RECT 99.635 51.56 99.915 52.32 ;
    RECT 99.635 50.8 99.915 51.56 ;
    RECT 99.635 50.04 99.915 50.8 ;
    RECT 99.635 49.28 99.915 50.04 ;
    RECT 99.635 48.52 99.915 49.28 ;
    RECT 99.635 47.76 99.915 48.52 ;
    RECT 99.635 11.28 99.915 12.04 ;
    RECT 99.635 47.0 99.915 47.76 ;
    RECT 99.635 46.24 99.915 47.0 ;
    RECT 99.635 45.48 99.915 46.24 ;
    RECT 99.635 44.72 99.915 45.48 ;
    RECT 99.635 43.96 99.915 44.72 ;
    RECT 99.635 43.2 99.915 43.96 ;
    RECT 99.635 42.44 99.915 43.2 ;
    RECT 99.635 41.68 99.915 42.44 ;
    RECT 99.635 40.92 99.915 41.68 ;
    RECT 99.635 40.16 99.915 40.92 ;
    RECT 99.635 109.3 99.915 110.77 ;
    RECT 99.635 39.4 99.915 40.16 ;
    RECT 99.635 38.64 99.915 39.4 ;
    RECT 99.635 37.88 99.915 38.64 ;
    RECT 99.635 37.12 99.915 37.88 ;
    RECT 99.635 36.36 99.915 37.12 ;
    RECT 99.635 35.6 99.915 36.36 ;
    RECT 99.635 34.84 99.915 35.6 ;
    RECT 99.635 34.08 99.915 34.84 ;
    RECT 99.635 107.78 99.915 108.54 ;
    RECT 99.635 33.32 99.915 34.08 ;
    RECT 99.635 107.02 99.915 107.78 ;
    RECT 99.635 32.56 99.915 33.32 ;
    RECT 99.635 106.26 99.915 107.02 ;
    RECT 99.635 105.5 99.915 106.26 ;
    RECT 99.635 104.74 99.915 105.5 ;
    RECT 99.635 103.98 99.915 104.74 ;
    RECT 99.635 103.22 99.915 103.98 ;
    RECT 99.635 102.46 99.915 103.22 ;
    RECT 99.635 101.7 99.915 102.46 ;
    RECT 99.635 100.94 99.915 101.7 ;
    RECT 96.535 31.8 96.815 32.56 ;
    RECT 96.535 31.04 96.815 31.8 ;
    RECT 96.535 30.28 96.815 31.04 ;
    RECT 96.535 29.52 96.815 30.28 ;
    RECT 96.535 28.76 96.815 29.52 ;
    RECT 96.535 28.0 96.815 28.76 ;
    RECT 96.535 27.24 96.815 28.0 ;
    RECT 96.535 26.48 96.815 27.24 ;
    RECT 96.535 100.18 96.815 100.94 ;
    RECT 96.535 25.72 96.815 26.48 ;
    RECT 96.535 99.42 96.815 100.18 ;
    RECT 96.535 24.96 96.815 25.72 ;
    RECT 96.535 98.66 96.815 99.42 ;
    RECT 96.535 97.9 96.815 98.66 ;
    RECT 96.535 97.14 96.815 97.9 ;
    RECT 96.535 96.38 96.815 97.14 ;
    RECT 96.535 95.62 96.815 96.38 ;
    RECT 96.535 94.86 96.815 95.62 ;
    RECT 96.535 94.1 96.815 94.86 ;
    RECT 96.535 93.34 96.815 94.1 ;
    RECT 96.535 24.2 96.815 24.96 ;
    RECT 96.535 23.44 96.815 24.2 ;
    RECT 96.535 22.68 96.815 23.44 ;
    RECT 96.535 21.92 96.815 22.68 ;
    RECT 96.535 21.16 96.815 21.92 ;
    RECT 96.535 20.4 96.815 21.16 ;
    RECT 96.535 19.64 96.815 20.4 ;
    RECT 96.535 18.88 96.815 19.64 ;
    RECT 96.535 92.58 96.815 93.34 ;
    RECT 96.535 18.12 96.815 18.88 ;
    RECT 96.535 91.82 96.815 92.58 ;
    RECT 96.535 17.36 96.815 18.12 ;
    RECT 96.535 91.06 96.815 91.82 ;
    RECT 96.535 90.3 96.815 91.06 ;
    RECT 96.535 89.54 96.815 90.3 ;
    RECT 96.535 88.78 96.815 89.54 ;
    RECT 96.535 88.02 96.815 88.78 ;
    RECT 96.535 87.26 96.815 88.02 ;
    RECT 96.535 86.5 96.815 87.26 ;
    RECT 96.535 85.74 96.815 86.5 ;
    RECT 96.535 84.98 96.815 85.74 ;
    RECT 96.535 84.22 96.815 84.98 ;
    RECT 96.535 83.46 96.815 84.22 ;
    RECT 96.535 82.7 96.815 83.46 ;
    RECT 96.535 81.94 96.815 82.7 ;
    RECT 96.535 81.18 96.815 81.94 ;
    RECT 96.535 80.42 96.815 81.18 ;
    RECT 96.535 79.66 96.815 80.42 ;
    RECT 96.535 78.9 96.815 79.66 ;
    RECT 96.535 78.14 96.815 78.9 ;
    RECT 96.535 77.38 96.815 78.14 ;
    RECT 96.535 76.62 96.815 77.38 ;
    RECT 96.535 75.86 96.815 76.62 ;
    RECT 96.535 75.1 96.815 75.86 ;
    RECT 96.535 74.34 96.815 75.1 ;
    RECT 96.535 73.58 96.815 74.34 ;
    RECT 96.535 72.82 96.815 73.58 ;
    RECT 96.535 72.06 96.815 72.82 ;
    RECT 96.535 71.3 96.815 72.06 ;
    RECT 96.535 70.54 96.815 71.3 ;
    RECT 96.535 69.78 96.815 70.54 ;
    RECT 96.535 69.02 96.815 69.78 ;
    RECT 96.535 68.26 96.815 69.02 ;
    RECT 96.535 67.5 96.815 68.26 ;
    RECT 96.535 66.74 96.815 67.5 ;
    RECT 96.535 65.98 96.815 66.74 ;
    RECT 96.535 65.22 96.815 65.98 ;
    RECT 96.535 64.46 96.815 65.22 ;
    RECT 96.535 63.7 96.815 64.46 ;
    RECT 96.535 62.94 96.815 63.7 ;
    RECT 96.535 108.54 96.815 109.3 ;
    RECT 96.535 62.18 96.815 62.94 ;
    RECT 96.535 61.42 96.815 62.18 ;
    RECT 96.535 60.66 96.815 61.42 ;
    RECT 96.535 59.92 96.815 60.66 ;
    RECT 96.535 59.16 96.815 59.92 ;
    RECT 96.535 58.4 96.815 59.16 ;
    RECT 96.535 57.64 96.815 58.4 ;
    RECT 96.535 56.88 96.815 57.64 ;
    RECT 96.535 56.12 96.815 56.88 ;
    RECT 96.535 55.36 96.815 56.12 ;
    RECT 96.535 16.6 96.815 17.36 ;
    RECT 96.535 15.84 96.815 16.6 ;
    RECT 96.535 15.08 96.815 15.84 ;
    RECT 96.535 14.32 96.815 15.08 ;
    RECT 96.535 13.56 96.815 14.32 ;
    RECT 96.535 12.8 96.815 13.56 ;
    RECT 96.535 12.04 96.815 12.8 ;
    RECT 96.535 9.81 96.815 11.28 ;
    RECT 96.535 54.6 96.815 55.36 ;
    RECT 96.535 53.84 96.815 54.6 ;
    RECT 96.535 53.08 96.815 53.84 ;
    RECT 96.535 52.32 96.815 53.08 ;
    RECT 96.535 51.56 96.815 52.32 ;
    RECT 96.535 50.8 96.815 51.56 ;
    RECT 96.535 50.04 96.815 50.8 ;
    RECT 96.535 49.28 96.815 50.04 ;
    RECT 96.535 48.52 96.815 49.28 ;
    RECT 96.535 47.76 96.815 48.52 ;
    RECT 96.535 11.28 96.815 12.04 ;
    RECT 96.535 47.0 96.815 47.76 ;
    RECT 96.535 46.24 96.815 47.0 ;
    RECT 96.535 45.48 96.815 46.24 ;
    RECT 96.535 44.72 96.815 45.48 ;
    RECT 96.535 43.96 96.815 44.72 ;
    RECT 96.535 43.2 96.815 43.96 ;
    RECT 96.535 42.44 96.815 43.2 ;
    RECT 96.535 41.68 96.815 42.44 ;
    RECT 96.535 40.92 96.815 41.68 ;
    RECT 96.535 40.16 96.815 40.92 ;
    RECT 96.535 109.3 96.815 110.77 ;
    RECT 96.535 39.4 96.815 40.16 ;
    RECT 96.535 38.64 96.815 39.4 ;
    RECT 96.535 37.88 96.815 38.64 ;
    RECT 96.535 37.12 96.815 37.88 ;
    RECT 96.535 36.36 96.815 37.12 ;
    RECT 96.535 35.6 96.815 36.36 ;
    RECT 96.535 34.84 96.815 35.6 ;
    RECT 96.535 34.08 96.815 34.84 ;
    RECT 96.535 107.78 96.815 108.54 ;
    RECT 96.535 33.32 96.815 34.08 ;
    RECT 96.535 107.02 96.815 107.78 ;
    RECT 96.535 32.56 96.815 33.32 ;
    RECT 96.535 106.26 96.815 107.02 ;
    RECT 96.535 105.5 96.815 106.26 ;
    RECT 96.535 104.74 96.815 105.5 ;
    RECT 96.535 103.98 96.815 104.74 ;
    RECT 96.535 103.22 96.815 103.98 ;
    RECT 96.535 102.46 96.815 103.22 ;
    RECT 96.535 101.7 96.815 102.46 ;
    RECT 96.535 100.94 96.815 101.7 ;
    RECT 93.435 31.8 93.715 32.56 ;
    RECT 93.435 31.04 93.715 31.8 ;
    RECT 93.435 30.28 93.715 31.04 ;
    RECT 93.435 29.52 93.715 30.28 ;
    RECT 93.435 28.76 93.715 29.52 ;
    RECT 93.435 28.0 93.715 28.76 ;
    RECT 93.435 27.24 93.715 28.0 ;
    RECT 93.435 26.48 93.715 27.24 ;
    RECT 93.435 100.18 93.715 100.94 ;
    RECT 93.435 25.72 93.715 26.48 ;
    RECT 93.435 99.42 93.715 100.18 ;
    RECT 93.435 24.96 93.715 25.72 ;
    RECT 93.435 98.66 93.715 99.42 ;
    RECT 93.435 97.9 93.715 98.66 ;
    RECT 93.435 97.14 93.715 97.9 ;
    RECT 93.435 96.38 93.715 97.14 ;
    RECT 93.435 95.62 93.715 96.38 ;
    RECT 93.435 94.86 93.715 95.62 ;
    RECT 93.435 94.1 93.715 94.86 ;
    RECT 93.435 93.34 93.715 94.1 ;
    RECT 93.435 24.2 93.715 24.96 ;
    RECT 93.435 23.44 93.715 24.2 ;
    RECT 93.435 22.68 93.715 23.44 ;
    RECT 93.435 21.92 93.715 22.68 ;
    RECT 93.435 21.16 93.715 21.92 ;
    RECT 93.435 20.4 93.715 21.16 ;
    RECT 93.435 19.64 93.715 20.4 ;
    RECT 93.435 18.88 93.715 19.64 ;
    RECT 93.435 92.58 93.715 93.34 ;
    RECT 93.435 18.12 93.715 18.88 ;
    RECT 93.435 91.82 93.715 92.58 ;
    RECT 93.435 17.36 93.715 18.12 ;
    RECT 93.435 91.06 93.715 91.82 ;
    RECT 93.435 90.3 93.715 91.06 ;
    RECT 93.435 89.54 93.715 90.3 ;
    RECT 93.435 88.78 93.715 89.54 ;
    RECT 93.435 88.02 93.715 88.78 ;
    RECT 93.435 87.26 93.715 88.02 ;
    RECT 93.435 86.5 93.715 87.26 ;
    RECT 93.435 85.74 93.715 86.5 ;
    RECT 93.435 84.98 93.715 85.74 ;
    RECT 93.435 84.22 93.715 84.98 ;
    RECT 93.435 83.46 93.715 84.22 ;
    RECT 93.435 82.7 93.715 83.46 ;
    RECT 93.435 81.94 93.715 82.7 ;
    RECT 93.435 81.18 93.715 81.94 ;
    RECT 93.435 80.42 93.715 81.18 ;
    RECT 93.435 79.66 93.715 80.42 ;
    RECT 93.435 78.9 93.715 79.66 ;
    RECT 93.435 78.14 93.715 78.9 ;
    RECT 93.435 77.38 93.715 78.14 ;
    RECT 93.435 76.62 93.715 77.38 ;
    RECT 93.435 75.86 93.715 76.62 ;
    RECT 93.435 75.1 93.715 75.86 ;
    RECT 93.435 74.34 93.715 75.1 ;
    RECT 93.435 73.58 93.715 74.34 ;
    RECT 93.435 72.82 93.715 73.58 ;
    RECT 93.435 72.06 93.715 72.82 ;
    RECT 93.435 71.3 93.715 72.06 ;
    RECT 93.435 70.54 93.715 71.3 ;
    RECT 93.435 69.78 93.715 70.54 ;
    RECT 93.435 69.02 93.715 69.78 ;
    RECT 93.435 68.26 93.715 69.02 ;
    RECT 93.435 67.5 93.715 68.26 ;
    RECT 93.435 66.74 93.715 67.5 ;
    RECT 93.435 65.98 93.715 66.74 ;
    RECT 93.435 65.22 93.715 65.98 ;
    RECT 93.435 64.46 93.715 65.22 ;
    RECT 93.435 63.7 93.715 64.46 ;
    RECT 93.435 62.94 93.715 63.7 ;
    RECT 93.435 108.54 93.715 109.3 ;
    RECT 93.435 62.18 93.715 62.94 ;
    RECT 93.435 61.42 93.715 62.18 ;
    RECT 93.435 60.66 93.715 61.42 ;
    RECT 93.435 59.92 93.715 60.66 ;
    RECT 93.435 59.16 93.715 59.92 ;
    RECT 93.435 58.4 93.715 59.16 ;
    RECT 93.435 57.64 93.715 58.4 ;
    RECT 93.435 56.88 93.715 57.64 ;
    RECT 93.435 56.12 93.715 56.88 ;
    RECT 93.435 55.36 93.715 56.12 ;
    RECT 93.435 16.6 93.715 17.36 ;
    RECT 93.435 15.84 93.715 16.6 ;
    RECT 93.435 15.08 93.715 15.84 ;
    RECT 93.435 14.32 93.715 15.08 ;
    RECT 93.435 13.56 93.715 14.32 ;
    RECT 93.435 12.8 93.715 13.56 ;
    RECT 93.435 12.04 93.715 12.8 ;
    RECT 93.435 9.81 93.715 11.28 ;
    RECT 93.435 54.6 93.715 55.36 ;
    RECT 93.435 53.84 93.715 54.6 ;
    RECT 93.435 53.08 93.715 53.84 ;
    RECT 93.435 52.32 93.715 53.08 ;
    RECT 93.435 51.56 93.715 52.32 ;
    RECT 93.435 50.8 93.715 51.56 ;
    RECT 93.435 50.04 93.715 50.8 ;
    RECT 93.435 49.28 93.715 50.04 ;
    RECT 93.435 48.52 93.715 49.28 ;
    RECT 93.435 47.76 93.715 48.52 ;
    RECT 93.435 11.28 93.715 12.04 ;
    RECT 93.435 47.0 93.715 47.76 ;
    RECT 93.435 46.24 93.715 47.0 ;
    RECT 93.435 45.48 93.715 46.24 ;
    RECT 93.435 44.72 93.715 45.48 ;
    RECT 93.435 43.96 93.715 44.72 ;
    RECT 93.435 43.2 93.715 43.96 ;
    RECT 93.435 42.44 93.715 43.2 ;
    RECT 93.435 41.68 93.715 42.44 ;
    RECT 93.435 40.92 93.715 41.68 ;
    RECT 93.435 40.16 93.715 40.92 ;
    RECT 93.435 109.3 93.715 110.77 ;
    RECT 93.435 39.4 93.715 40.16 ;
    RECT 93.435 38.64 93.715 39.4 ;
    RECT 93.435 37.88 93.715 38.64 ;
    RECT 93.435 37.12 93.715 37.88 ;
    RECT 93.435 36.36 93.715 37.12 ;
    RECT 93.435 35.6 93.715 36.36 ;
    RECT 93.435 34.84 93.715 35.6 ;
    RECT 93.435 34.08 93.715 34.84 ;
    RECT 93.435 107.78 93.715 108.54 ;
    RECT 93.435 33.32 93.715 34.08 ;
    RECT 93.435 107.02 93.715 107.78 ;
    RECT 93.435 32.56 93.715 33.32 ;
    RECT 93.435 106.26 93.715 107.02 ;
    RECT 93.435 105.5 93.715 106.26 ;
    RECT 93.435 104.74 93.715 105.5 ;
    RECT 93.435 103.98 93.715 104.74 ;
    RECT 93.435 103.22 93.715 103.98 ;
    RECT 93.435 102.46 93.715 103.22 ;
    RECT 93.435 101.7 93.715 102.46 ;
    RECT 93.435 100.94 93.715 101.7 ;
    RECT 105.835 31.8 106.115 32.56 ;
    RECT 105.835 31.04 106.115 31.8 ;
    RECT 105.835 30.28 106.115 31.04 ;
    RECT 105.835 29.52 106.115 30.28 ;
    RECT 105.835 28.76 106.115 29.52 ;
    RECT 105.835 28.0 106.115 28.76 ;
    RECT 105.835 27.24 106.115 28.0 ;
    RECT 105.835 26.48 106.115 27.24 ;
    RECT 105.835 100.18 106.115 100.94 ;
    RECT 105.835 25.72 106.115 26.48 ;
    RECT 105.835 99.42 106.115 100.18 ;
    RECT 105.835 24.96 106.115 25.72 ;
    RECT 105.835 98.66 106.115 99.42 ;
    RECT 105.835 97.9 106.115 98.66 ;
    RECT 105.835 97.14 106.115 97.9 ;
    RECT 105.835 96.38 106.115 97.14 ;
    RECT 105.835 95.62 106.115 96.38 ;
    RECT 105.835 94.86 106.115 95.62 ;
    RECT 105.835 94.1 106.115 94.86 ;
    RECT 105.835 93.34 106.115 94.1 ;
    RECT 105.835 24.2 106.115 24.96 ;
    RECT 105.835 23.44 106.115 24.2 ;
    RECT 105.835 22.68 106.115 23.44 ;
    RECT 105.835 21.92 106.115 22.68 ;
    RECT 105.835 21.16 106.115 21.92 ;
    RECT 105.835 20.4 106.115 21.16 ;
    RECT 105.835 19.64 106.115 20.4 ;
    RECT 105.835 18.88 106.115 19.64 ;
    RECT 105.835 92.58 106.115 93.34 ;
    RECT 105.835 18.12 106.115 18.88 ;
    RECT 105.835 91.82 106.115 92.58 ;
    RECT 105.835 17.36 106.115 18.12 ;
    RECT 105.835 91.06 106.115 91.82 ;
    RECT 105.835 90.3 106.115 91.06 ;
    RECT 105.835 89.54 106.115 90.3 ;
    RECT 105.835 88.78 106.115 89.54 ;
    RECT 105.835 88.02 106.115 88.78 ;
    RECT 105.835 87.26 106.115 88.02 ;
    RECT 105.835 86.5 106.115 87.26 ;
    RECT 105.835 85.74 106.115 86.5 ;
    RECT 105.835 84.98 106.115 85.74 ;
    RECT 105.835 84.22 106.115 84.98 ;
    RECT 105.835 83.46 106.115 84.22 ;
    RECT 105.835 82.7 106.115 83.46 ;
    RECT 105.835 81.94 106.115 82.7 ;
    RECT 105.835 81.18 106.115 81.94 ;
    RECT 105.835 80.42 106.115 81.18 ;
    RECT 105.835 79.66 106.115 80.42 ;
    RECT 105.835 78.9 106.115 79.66 ;
    RECT 105.835 78.14 106.115 78.9 ;
    RECT 105.835 77.38 106.115 78.14 ;
    RECT 105.835 76.62 106.115 77.38 ;
    RECT 105.835 75.86 106.115 76.62 ;
    RECT 105.835 75.1 106.115 75.86 ;
    RECT 105.835 74.34 106.115 75.1 ;
    RECT 105.835 73.58 106.115 74.34 ;
    RECT 105.835 72.82 106.115 73.58 ;
    RECT 105.835 72.06 106.115 72.82 ;
    RECT 105.835 71.3 106.115 72.06 ;
    RECT 105.835 70.54 106.115 71.3 ;
    RECT 105.835 69.78 106.115 70.54 ;
    RECT 105.835 69.02 106.115 69.78 ;
    RECT 105.835 68.26 106.115 69.02 ;
    RECT 105.835 67.5 106.115 68.26 ;
    RECT 105.835 66.74 106.115 67.5 ;
    RECT 105.835 65.98 106.115 66.74 ;
    RECT 105.835 65.22 106.115 65.98 ;
    RECT 105.835 64.46 106.115 65.22 ;
    RECT 105.835 63.7 106.115 64.46 ;
    RECT 105.835 62.94 106.115 63.7 ;
    RECT 105.835 108.54 106.115 109.3 ;
    RECT 105.835 62.18 106.115 62.94 ;
    RECT 105.835 61.42 106.115 62.18 ;
    RECT 105.835 60.66 106.115 61.42 ;
    RECT 105.835 59.92 106.115 60.66 ;
    RECT 105.835 59.16 106.115 59.92 ;
    RECT 105.835 58.4 106.115 59.16 ;
    RECT 105.835 57.64 106.115 58.4 ;
    RECT 105.835 56.88 106.115 57.64 ;
    RECT 105.835 56.12 106.115 56.88 ;
    RECT 105.835 55.36 106.115 56.12 ;
    RECT 105.835 16.6 106.115 17.36 ;
    RECT 105.835 15.84 106.115 16.6 ;
    RECT 105.835 15.08 106.115 15.84 ;
    RECT 105.835 14.32 106.115 15.08 ;
    RECT 105.835 13.56 106.115 14.32 ;
    RECT 105.835 12.8 106.115 13.56 ;
    RECT 105.835 12.04 106.115 12.8 ;
    RECT 105.835 9.81 106.115 11.28 ;
    RECT 105.835 54.6 106.115 55.36 ;
    RECT 105.835 53.84 106.115 54.6 ;
    RECT 105.835 53.08 106.115 53.84 ;
    RECT 105.835 52.32 106.115 53.08 ;
    RECT 105.835 51.56 106.115 52.32 ;
    RECT 105.835 50.8 106.115 51.56 ;
    RECT 105.835 50.04 106.115 50.8 ;
    RECT 105.835 49.28 106.115 50.04 ;
    RECT 105.835 48.52 106.115 49.28 ;
    RECT 105.835 47.76 106.115 48.52 ;
    RECT 105.835 11.28 106.115 12.04 ;
    RECT 105.835 47.0 106.115 47.76 ;
    RECT 105.835 46.24 106.115 47.0 ;
    RECT 105.835 45.48 106.115 46.24 ;
    RECT 105.835 44.72 106.115 45.48 ;
    RECT 105.835 43.96 106.115 44.72 ;
    RECT 105.835 43.2 106.115 43.96 ;
    RECT 105.835 42.44 106.115 43.2 ;
    RECT 105.835 41.68 106.115 42.44 ;
    RECT 105.835 40.92 106.115 41.68 ;
    RECT 105.835 40.16 106.115 40.92 ;
    RECT 105.835 109.3 106.115 110.77 ;
    RECT 105.835 39.4 106.115 40.16 ;
    RECT 105.835 38.64 106.115 39.4 ;
    RECT 105.835 37.88 106.115 38.64 ;
    RECT 105.835 37.12 106.115 37.88 ;
    RECT 105.835 36.36 106.115 37.12 ;
    RECT 105.835 35.6 106.115 36.36 ;
    RECT 105.835 34.84 106.115 35.6 ;
    RECT 105.835 34.08 106.115 34.84 ;
    RECT 105.835 107.78 106.115 108.54 ;
    RECT 105.835 33.32 106.115 34.08 ;
    RECT 105.835 107.02 106.115 107.78 ;
    RECT 105.835 32.56 106.115 33.32 ;
    RECT 105.835 106.26 106.115 107.02 ;
    RECT 105.835 105.5 106.115 106.26 ;
    RECT 105.835 104.74 106.115 105.5 ;
    RECT 105.835 103.98 106.115 104.74 ;
    RECT 105.835 103.22 106.115 103.98 ;
    RECT 105.835 102.46 106.115 103.22 ;
    RECT 105.835 101.7 106.115 102.46 ;
    RECT 105.835 100.94 106.115 101.7 ;
    RECT 87.235 31.8 87.515 32.56 ;
    RECT 87.235 31.04 87.515 31.8 ;
    RECT 87.235 30.28 87.515 31.04 ;
    RECT 87.235 29.52 87.515 30.28 ;
    RECT 87.235 28.76 87.515 29.52 ;
    RECT 87.235 28.0 87.515 28.76 ;
    RECT 87.235 27.24 87.515 28.0 ;
    RECT 87.235 26.48 87.515 27.24 ;
    RECT 87.235 100.18 87.515 100.94 ;
    RECT 87.235 25.72 87.515 26.48 ;
    RECT 87.235 99.42 87.515 100.18 ;
    RECT 87.235 24.96 87.515 25.72 ;
    RECT 87.235 98.66 87.515 99.42 ;
    RECT 87.235 97.9 87.515 98.66 ;
    RECT 87.235 97.14 87.515 97.9 ;
    RECT 87.235 96.38 87.515 97.14 ;
    RECT 87.235 95.62 87.515 96.38 ;
    RECT 87.235 94.86 87.515 95.62 ;
    RECT 87.235 94.1 87.515 94.86 ;
    RECT 87.235 93.34 87.515 94.1 ;
    RECT 87.235 24.2 87.515 24.96 ;
    RECT 87.235 23.44 87.515 24.2 ;
    RECT 87.235 22.68 87.515 23.44 ;
    RECT 87.235 21.92 87.515 22.68 ;
    RECT 87.235 21.16 87.515 21.92 ;
    RECT 87.235 20.4 87.515 21.16 ;
    RECT 87.235 19.64 87.515 20.4 ;
    RECT 87.235 18.88 87.515 19.64 ;
    RECT 87.235 92.58 87.515 93.34 ;
    RECT 87.235 18.12 87.515 18.88 ;
    RECT 87.235 91.82 87.515 92.58 ;
    RECT 87.235 17.36 87.515 18.12 ;
    RECT 87.235 91.06 87.515 91.82 ;
    RECT 87.235 90.3 87.515 91.06 ;
    RECT 87.235 89.54 87.515 90.3 ;
    RECT 87.235 88.78 87.515 89.54 ;
    RECT 87.235 88.02 87.515 88.78 ;
    RECT 87.235 87.26 87.515 88.02 ;
    RECT 87.235 86.5 87.515 87.26 ;
    RECT 87.235 85.74 87.515 86.5 ;
    RECT 87.235 84.98 87.515 85.74 ;
    RECT 87.235 84.22 87.515 84.98 ;
    RECT 87.235 83.46 87.515 84.22 ;
    RECT 87.235 82.7 87.515 83.46 ;
    RECT 87.235 81.94 87.515 82.7 ;
    RECT 87.235 81.18 87.515 81.94 ;
    RECT 87.235 80.42 87.515 81.18 ;
    RECT 87.235 79.66 87.515 80.42 ;
    RECT 87.235 78.9 87.515 79.66 ;
    RECT 87.235 78.14 87.515 78.9 ;
    RECT 87.235 77.38 87.515 78.14 ;
    RECT 87.235 76.62 87.515 77.38 ;
    RECT 87.235 75.86 87.515 76.62 ;
    RECT 87.235 75.1 87.515 75.86 ;
    RECT 87.235 74.34 87.515 75.1 ;
    RECT 87.235 73.58 87.515 74.34 ;
    RECT 87.235 72.82 87.515 73.58 ;
    RECT 87.235 72.06 87.515 72.82 ;
    RECT 87.235 71.3 87.515 72.06 ;
    RECT 87.235 70.54 87.515 71.3 ;
    RECT 87.235 69.78 87.515 70.54 ;
    RECT 87.235 69.02 87.515 69.78 ;
    RECT 87.235 68.26 87.515 69.02 ;
    RECT 87.235 67.5 87.515 68.26 ;
    RECT 87.235 66.74 87.515 67.5 ;
    RECT 87.235 65.98 87.515 66.74 ;
    RECT 87.235 65.22 87.515 65.98 ;
    RECT 87.235 64.46 87.515 65.22 ;
    RECT 87.235 63.7 87.515 64.46 ;
    RECT 87.235 62.94 87.515 63.7 ;
    RECT 87.235 108.54 87.515 109.3 ;
    RECT 87.235 62.18 87.515 62.94 ;
    RECT 87.235 61.42 87.515 62.18 ;
    RECT 87.235 60.66 87.515 61.42 ;
    RECT 87.235 59.92 87.515 60.66 ;
    RECT 87.235 59.16 87.515 59.92 ;
    RECT 87.235 58.4 87.515 59.16 ;
    RECT 87.235 57.64 87.515 58.4 ;
    RECT 87.235 56.88 87.515 57.64 ;
    RECT 87.235 56.12 87.515 56.88 ;
    RECT 87.235 55.36 87.515 56.12 ;
    RECT 87.235 16.6 87.515 17.36 ;
    RECT 87.235 15.84 87.515 16.6 ;
    RECT 87.235 15.08 87.515 15.84 ;
    RECT 87.235 14.32 87.515 15.08 ;
    RECT 87.235 13.56 87.515 14.32 ;
    RECT 87.235 12.8 87.515 13.56 ;
    RECT 87.235 12.04 87.515 12.8 ;
    RECT 87.235 9.81 87.515 11.28 ;
    RECT 87.235 54.6 87.515 55.36 ;
    RECT 87.235 53.84 87.515 54.6 ;
    RECT 87.235 53.08 87.515 53.84 ;
    RECT 87.235 52.32 87.515 53.08 ;
    RECT 87.235 51.56 87.515 52.32 ;
    RECT 87.235 50.8 87.515 51.56 ;
    RECT 87.235 50.04 87.515 50.8 ;
    RECT 87.235 49.28 87.515 50.04 ;
    RECT 87.235 48.52 87.515 49.28 ;
    RECT 87.235 47.76 87.515 48.52 ;
    RECT 87.235 11.28 87.515 12.04 ;
    RECT 87.235 47.0 87.515 47.76 ;
    RECT 87.235 46.24 87.515 47.0 ;
    RECT 87.235 45.48 87.515 46.24 ;
    RECT 87.235 44.72 87.515 45.48 ;
    RECT 87.235 43.96 87.515 44.72 ;
    RECT 87.235 43.2 87.515 43.96 ;
    RECT 87.235 42.44 87.515 43.2 ;
    RECT 87.235 41.68 87.515 42.44 ;
    RECT 87.235 40.92 87.515 41.68 ;
    RECT 87.235 40.16 87.515 40.92 ;
    RECT 87.235 109.3 87.515 110.77 ;
    RECT 87.235 39.4 87.515 40.16 ;
    RECT 87.235 38.64 87.515 39.4 ;
    RECT 87.235 37.88 87.515 38.64 ;
    RECT 87.235 37.12 87.515 37.88 ;
    RECT 87.235 36.36 87.515 37.12 ;
    RECT 87.235 35.6 87.515 36.36 ;
    RECT 87.235 34.84 87.515 35.6 ;
    RECT 87.235 34.08 87.515 34.84 ;
    RECT 87.235 107.78 87.515 108.54 ;
    RECT 87.235 33.32 87.515 34.08 ;
    RECT 87.235 107.02 87.515 107.78 ;
    RECT 87.235 32.56 87.515 33.32 ;
    RECT 87.235 106.26 87.515 107.02 ;
    RECT 87.235 105.5 87.515 106.26 ;
    RECT 87.235 104.74 87.515 105.5 ;
    RECT 87.235 103.98 87.515 104.74 ;
    RECT 87.235 103.22 87.515 103.98 ;
    RECT 87.235 102.46 87.515 103.22 ;
    RECT 87.235 101.7 87.515 102.46 ;
    RECT 87.235 100.94 87.515 101.7 ;
    RECT 108.935 31.8 109.215 32.56 ;
    RECT 108.935 31.04 109.215 31.8 ;
    RECT 108.935 30.28 109.215 31.04 ;
    RECT 108.935 29.52 109.215 30.28 ;
    RECT 108.935 28.76 109.215 29.52 ;
    RECT 108.935 28.0 109.215 28.76 ;
    RECT 108.935 27.24 109.215 28.0 ;
    RECT 108.935 26.48 109.215 27.24 ;
    RECT 108.935 100.18 109.215 100.94 ;
    RECT 108.935 25.72 109.215 26.48 ;
    RECT 108.935 99.42 109.215 100.18 ;
    RECT 108.935 24.96 109.215 25.72 ;
    RECT 108.935 98.66 109.215 99.42 ;
    RECT 108.935 97.9 109.215 98.66 ;
    RECT 108.935 97.14 109.215 97.9 ;
    RECT 108.935 96.38 109.215 97.14 ;
    RECT 108.935 95.62 109.215 96.38 ;
    RECT 108.935 94.86 109.215 95.62 ;
    RECT 108.935 94.1 109.215 94.86 ;
    RECT 108.935 93.34 109.215 94.1 ;
    RECT 108.935 24.2 109.215 24.96 ;
    RECT 108.935 23.44 109.215 24.2 ;
    RECT 108.935 22.68 109.215 23.44 ;
    RECT 108.935 21.92 109.215 22.68 ;
    RECT 108.935 21.16 109.215 21.92 ;
    RECT 108.935 20.4 109.215 21.16 ;
    RECT 108.935 19.64 109.215 20.4 ;
    RECT 108.935 18.88 109.215 19.64 ;
    RECT 108.935 92.58 109.215 93.34 ;
    RECT 108.935 18.12 109.215 18.88 ;
    RECT 108.935 91.82 109.215 92.58 ;
    RECT 108.935 17.36 109.215 18.12 ;
    RECT 108.935 91.06 109.215 91.82 ;
    RECT 108.935 90.3 109.215 91.06 ;
    RECT 108.935 89.54 109.215 90.3 ;
    RECT 108.935 88.78 109.215 89.54 ;
    RECT 108.935 88.02 109.215 88.78 ;
    RECT 108.935 87.26 109.215 88.02 ;
    RECT 108.935 86.5 109.215 87.26 ;
    RECT 108.935 85.74 109.215 86.5 ;
    RECT 108.935 84.98 109.215 85.74 ;
    RECT 108.935 84.22 109.215 84.98 ;
    RECT 108.935 83.46 109.215 84.22 ;
    RECT 108.935 82.7 109.215 83.46 ;
    RECT 108.935 81.94 109.215 82.7 ;
    RECT 108.935 81.18 109.215 81.94 ;
    RECT 108.935 80.42 109.215 81.18 ;
    RECT 108.935 79.66 109.215 80.42 ;
    RECT 108.935 78.9 109.215 79.66 ;
    RECT 108.935 78.14 109.215 78.9 ;
    RECT 108.935 77.38 109.215 78.14 ;
    RECT 108.935 76.62 109.215 77.38 ;
    RECT 108.935 75.86 109.215 76.62 ;
    RECT 108.935 75.1 109.215 75.86 ;
    RECT 108.935 74.34 109.215 75.1 ;
    RECT 108.935 73.58 109.215 74.34 ;
    RECT 108.935 72.82 109.215 73.58 ;
    RECT 108.935 72.06 109.215 72.82 ;
    RECT 108.935 71.3 109.215 72.06 ;
    RECT 108.935 70.54 109.215 71.3 ;
    RECT 108.935 69.78 109.215 70.54 ;
    RECT 108.935 69.02 109.215 69.78 ;
    RECT 108.935 68.26 109.215 69.02 ;
    RECT 108.935 67.5 109.215 68.26 ;
    RECT 108.935 66.74 109.215 67.5 ;
    RECT 108.935 65.98 109.215 66.74 ;
    RECT 108.935 65.22 109.215 65.98 ;
    RECT 108.935 64.46 109.215 65.22 ;
    RECT 108.935 63.7 109.215 64.46 ;
    RECT 108.935 62.94 109.215 63.7 ;
    RECT 108.935 108.54 109.215 109.3 ;
    RECT 108.935 62.18 109.215 62.94 ;
    RECT 108.935 61.42 109.215 62.18 ;
    RECT 108.935 60.66 109.215 61.42 ;
    RECT 108.935 59.92 109.215 60.66 ;
    RECT 108.935 59.16 109.215 59.92 ;
    RECT 108.935 58.4 109.215 59.16 ;
    RECT 108.935 57.64 109.215 58.4 ;
    RECT 108.935 56.88 109.215 57.64 ;
    RECT 108.935 56.12 109.215 56.88 ;
    RECT 108.935 55.36 109.215 56.12 ;
    RECT 108.935 16.6 109.215 17.36 ;
    RECT 108.935 15.84 109.215 16.6 ;
    RECT 108.935 15.08 109.215 15.84 ;
    RECT 108.935 14.32 109.215 15.08 ;
    RECT 108.935 13.56 109.215 14.32 ;
    RECT 108.935 12.8 109.215 13.56 ;
    RECT 108.935 12.04 109.215 12.8 ;
    RECT 108.935 9.81 109.215 11.28 ;
    RECT 108.935 54.6 109.215 55.36 ;
    RECT 108.935 53.84 109.215 54.6 ;
    RECT 108.935 53.08 109.215 53.84 ;
    RECT 108.935 52.32 109.215 53.08 ;
    RECT 108.935 51.56 109.215 52.32 ;
    RECT 108.935 50.8 109.215 51.56 ;
    RECT 108.935 50.04 109.215 50.8 ;
    RECT 108.935 49.28 109.215 50.04 ;
    RECT 108.935 48.52 109.215 49.28 ;
    RECT 108.935 47.76 109.215 48.52 ;
    RECT 108.935 11.28 109.215 12.04 ;
    RECT 108.935 47.0 109.215 47.76 ;
    RECT 108.935 46.24 109.215 47.0 ;
    RECT 108.935 45.48 109.215 46.24 ;
    RECT 108.935 44.72 109.215 45.48 ;
    RECT 108.935 43.96 109.215 44.72 ;
    RECT 108.935 43.2 109.215 43.96 ;
    RECT 108.935 42.44 109.215 43.2 ;
    RECT 108.935 41.68 109.215 42.44 ;
    RECT 108.935 40.92 109.215 41.68 ;
    RECT 108.935 40.16 109.215 40.92 ;
    RECT 108.935 109.3 109.215 110.77 ;
    RECT 108.935 39.4 109.215 40.16 ;
    RECT 108.935 38.64 109.215 39.4 ;
    RECT 108.935 37.88 109.215 38.64 ;
    RECT 108.935 37.12 109.215 37.88 ;
    RECT 108.935 36.36 109.215 37.12 ;
    RECT 108.935 35.6 109.215 36.36 ;
    RECT 108.935 34.84 109.215 35.6 ;
    RECT 108.935 34.08 109.215 34.84 ;
    RECT 108.935 107.78 109.215 108.54 ;
    RECT 108.935 33.32 109.215 34.08 ;
    RECT 108.935 107.02 109.215 107.78 ;
    RECT 108.935 32.56 109.215 33.32 ;
    RECT 108.935 106.26 109.215 107.02 ;
    RECT 108.935 105.5 109.215 106.26 ;
    RECT 108.935 104.74 109.215 105.5 ;
    RECT 108.935 103.98 109.215 104.74 ;
    RECT 108.935 103.22 109.215 103.98 ;
    RECT 108.935 102.46 109.215 103.22 ;
    RECT 108.935 101.7 109.215 102.46 ;
    RECT 108.935 100.94 109.215 101.7 ;
    RECT 26.78 110.77 27.32 111.115 ;
    RECT 27.8 110.77 28.02 111.115 ;
    RECT 28.5 110.77 28.72 111.115 ;
    RECT 29.2 110.77 30.815 111.115 ;
    RECT 31.295 110.77 31.515 111.115 ;
    RECT 31.995 110.77 32.21 111.115 ;
    RECT 32.69 110.77 32.91 111.115 ;
    RECT 33.39 110.77 33.61 111.115 ;
    RECT 34.09 110.77 34.31 111.115 ;
    RECT 34.79 110.77 35.005 111.115 ;
    RECT 35.485 110.77 36.405 111.115 ;
    RECT 36.885 110.77 37.105 111.115 ;
    RECT 37.585 110.77 37.8 111.115 ;
    RECT 38.28 110.77 38.5 111.115 ;
    RECT 38.98 110.77 39.2 111.115 ;
    RECT 39.68 110.77 39.895 111.115 ;
    RECT 40.375 110.77 40.595 111.115 ;
    RECT 41.075 110.77 41.995 111.115 ;
    RECT 42.475 110.77 42.69 111.115 ;
    RECT 43.17 110.77 43.39 111.115 ;
    RECT 43.87 110.77 44.09 111.115 ;
    RECT 44.57 110.77 44.79 111.115 ;
    RECT 45.27 110.77 45.485 111.115 ;
    RECT 45.965 110.77 46.185 111.115 ;
    RECT 46.665 110.77 47.58 111.115 ;
    RECT 48.06 110.77 48.28 111.115 ;
    RECT 48.76 110.77 48.98 111.115 ;
    RECT 49.46 110.77 49.68 111.115 ;
    RECT 50.16 110.77 50.375 111.115 ;
    RECT 50.855 110.77 51.775 111.115 ;
    RECT 52.255 110.77 53.17 111.115 ;
    RECT 53.65 110.77 53.87 111.115 ;
    RECT 54.35 110.77 54.57 111.115 ;
    RECT 55.05 110.77 55.265 111.115 ;
    RECT 55.745 110.77 55.965 111.115 ;
    RECT 56.445 110.77 56.665 111.115 ;
    RECT 57.145 110.77 58.06 111.115 ;
    RECT 58.54 110.77 59.46 111.115 ;
    RECT 59.94 110.77 60.16 111.115 ;
    RECT 60.64 110.77 60.855 111.115 ;
    RECT 61.335 110.77 61.555 111.115 ;
    RECT 62.035 110.77 62.25 111.115 ;
    RECT 62.73 110.77 63.65 111.115 ;
    RECT 64.13 110.77 64.345 111.115 ;
    RECT 64.825 110.77 65.045 111.115 ;
    RECT 65.525 110.77 65.745 111.115 ;
    RECT 66.225 110.77 66.445 111.115 ;
    RECT 66.925 110.77 67.14 111.115 ;
    RECT 67.62 110.77 67.84 111.115 ;
    RECT 68.32 110.77 69.235 111.115 ;
    RECT 69.715 110.77 69.935 111.115 ;
    RECT 70.415 110.77 70.635 111.115 ;
    RECT 71.115 110.77 71.335 111.115 ;
    RECT 71.815 110.77 72.035 111.115 ;
    RECT 72.515 110.77 72.735 111.115 ;
    RECT 73.215 110.77 73.435 111.115 ;
    RECT 73.915 110.77 74.835 111.115 ;
    RECT 75.315 110.77 75.535 111.115 ;
    RECT 77.4 110.77 77.62 111.115 ;
    RECT 78.1 110.77 78.32 111.115 ;
    RECT 78.8 110.77 79.02 111.115 ;
    RECT 79.5 110.77 80.515 111.115 ;
    RECT 80.515 110.605 80.795 111.115 ;
    RECT 80.795 110.77 81.115 111.115 ;
    RECT 81.595 110.77 81.815 111.115 ;
    RECT 82.295 110.77 82.515 111.115 ;
    RECT 82.995 110.77 83.055 111.115 ;
    RECT 83.055 110.605 83.335 111.115 ;
    RECT 83.335 110.77 83.435 111.115 ;
    RECT 26.71 9.81 26.88 23.44 ;
    RECT 26.88 9.81 27.16 23.53 ;
    RECT 27.16 9.81 27.32 23.44 ;
    RECT 27.8 9.81 28.02 23.44 ;
    RECT 28.5 9.81 28.72 23.44 ;
    RECT 29.2 9.81 30.815 23.44 ;
    RECT 31.295 9.81 31.515 23.44 ;
    RECT 31.995 9.81 32.21 23.44 ;
    RECT 32.69 9.81 32.91 23.44 ;
    RECT 33.39 9.81 33.61 23.44 ;
    RECT 34.09 9.81 34.31 23.44 ;
    RECT 34.79 9.81 35.005 23.44 ;
    RECT 35.485 9.81 36.405 23.44 ;
    RECT 36.885 9.81 37.105 23.44 ;
    RECT 37.585 9.81 37.8 23.44 ;
    RECT 38.28 9.81 38.5 23.44 ;
    RECT 38.98 9.81 39.2 23.44 ;
    RECT 39.68 9.81 39.895 23.44 ;
    RECT 40.375 9.81 40.595 23.44 ;
    RECT 41.075 9.81 41.995 23.44 ;
    RECT 42.475 9.81 42.69 23.44 ;
    RECT 43.17 9.81 43.39 23.44 ;
    RECT 43.87 9.81 44.09 23.44 ;
    RECT 44.57 9.81 44.79 23.44 ;
    RECT 45.27 9.81 45.485 23.44 ;
    RECT 45.965 9.81 46.185 23.44 ;
    RECT 46.665 9.81 47.58 23.44 ;
    RECT 48.06 9.81 48.28 23.44 ;
    RECT 48.76 9.81 48.98 23.44 ;
    RECT 49.46 9.81 49.68 23.44 ;
    RECT 50.16 9.81 50.375 23.44 ;
    RECT 50.855 9.81 51.775 23.44 ;
    RECT 52.255 9.81 53.17 23.44 ;
    RECT 53.65 9.81 53.87 23.44 ;
    RECT 54.35 9.81 54.57 23.44 ;
    RECT 55.05 9.81 55.265 23.44 ;
    RECT 55.745 9.81 55.965 23.44 ;
    RECT 56.445 9.81 56.665 23.44 ;
    RECT 57.145 9.81 58.06 23.44 ;
    RECT 58.54 9.81 59.46 23.44 ;
    RECT 59.94 9.81 60.16 23.44 ;
    RECT 60.64 9.81 60.855 23.44 ;
    RECT 61.335 9.81 61.555 23.44 ;
    RECT 62.035 9.81 62.25 23.44 ;
    RECT 62.73 9.81 63.65 23.44 ;
    RECT 64.13 9.81 64.345 23.44 ;
    RECT 64.825 9.81 65.045 23.44 ;
    RECT 65.525 9.81 65.745 23.44 ;
    RECT 66.225 9.81 66.445 23.44 ;
    RECT 66.925 9.81 67.14 23.44 ;
    RECT 67.62 9.81 67.84 23.44 ;
    RECT 68.32 9.81 69.235 23.44 ;
    RECT 69.715 9.81 69.935 23.44 ;
    RECT 70.415 9.81 70.635 23.44 ;
    RECT 71.115 9.81 71.335 23.44 ;
    RECT 71.815 9.81 72.035 23.44 ;
    RECT 72.515 9.81 72.735 23.44 ;
    RECT 73.215 9.81 73.435 23.44 ;
    RECT 73.915 9.81 74.835 23.44 ;
    RECT 75.315 9.81 75.535 23.44 ;
    RECT 76.015 9.81 76.225 23.44 ;
    RECT 76.705 9.81 76.92 23.44 ;
    RECT 77.4 9.81 77.62 23.44 ;
    RECT 78.1 9.81 78.32 23.44 ;
    RECT 78.8 9.81 79.02 23.44 ;
    RECT 79.5 9.81 81.115 23.44 ;
    RECT 81.595 9.81 81.815 23.44 ;
    RECT 82.295 9.81 82.515 23.44 ;
    RECT 82.995 9.81 83.055 23.44 ;
    RECT 83.055 9.81 83.335 23.53 ;
    RECT 83.335 9.81 83.505 23.44 ;
    RECT 26.71 107.78 26.88 108.54 ;
    RECT 26.88 107.69 27.16 108.63 ;
    RECT 27.16 107.78 27.32 108.54 ;
    RECT 27.8 107.78 28.02 108.54 ;
    RECT 28.5 107.78 28.72 108.54 ;
    RECT 29.2 107.78 30.815 108.54 ;
    RECT 31.295 107.78 31.515 108.54 ;
    RECT 31.995 107.78 32.21 108.54 ;
    RECT 32.69 107.78 32.91 108.54 ;
    RECT 33.39 107.78 33.61 108.54 ;
    RECT 34.09 107.78 34.31 108.54 ;
    RECT 34.79 107.78 35.005 108.54 ;
    RECT 35.485 107.78 36.405 108.54 ;
    RECT 36.885 107.78 37.105 108.54 ;
    RECT 37.585 107.78 37.8 108.54 ;
    RECT 38.28 107.78 38.5 108.54 ;
    RECT 38.98 107.78 39.2 108.54 ;
    RECT 39.68 107.78 39.895 108.54 ;
    RECT 40.375 107.78 40.595 108.54 ;
    RECT 41.075 107.78 41.995 108.54 ;
    RECT 42.475 107.78 42.69 108.54 ;
    RECT 43.17 107.78 43.39 108.54 ;
    RECT 43.87 107.78 44.09 108.54 ;
    RECT 44.57 107.78 44.79 108.54 ;
    RECT 45.27 107.78 45.485 108.54 ;
    RECT 45.965 107.78 46.185 108.54 ;
    RECT 46.665 107.78 47.58 108.54 ;
    RECT 48.06 107.78 48.28 108.54 ;
    RECT 48.76 107.78 48.98 108.54 ;
    RECT 49.46 107.78 49.68 108.54 ;
    RECT 50.16 107.78 50.375 108.54 ;
    RECT 50.855 107.78 51.775 108.54 ;
    RECT 52.255 107.78 53.17 108.54 ;
    RECT 53.65 107.78 53.87 108.54 ;
    RECT 54.35 107.78 54.57 108.54 ;
    RECT 55.05 107.78 55.265 108.54 ;
    RECT 55.745 107.78 55.965 108.54 ;
    RECT 56.445 107.78 56.665 108.54 ;
    RECT 57.145 107.78 58.06 108.54 ;
    RECT 58.54 107.78 59.46 108.54 ;
    RECT 59.94 107.78 60.16 108.54 ;
    RECT 60.64 107.78 60.855 108.54 ;
    RECT 61.335 107.78 61.555 108.54 ;
    RECT 62.035 107.78 62.25 108.54 ;
    RECT 62.73 107.78 63.65 108.54 ;
    RECT 64.13 107.78 64.345 108.54 ;
    RECT 64.825 107.78 65.045 108.54 ;
    RECT 65.525 107.78 65.745 108.54 ;
    RECT 66.225 107.78 66.445 108.54 ;
    RECT 66.925 107.78 67.14 108.54 ;
    RECT 67.62 107.78 67.84 108.54 ;
    RECT 68.32 107.78 69.235 108.54 ;
    RECT 69.715 107.78 69.935 108.54 ;
    RECT 70.415 107.78 70.635 108.54 ;
    RECT 71.115 107.78 71.335 108.54 ;
    RECT 71.815 107.78 72.035 108.54 ;
    RECT 72.515 107.78 72.735 108.54 ;
    RECT 73.215 107.78 73.435 108.54 ;
    RECT 73.915 107.78 74.835 108.54 ;
    RECT 75.315 107.78 75.535 108.54 ;
    RECT 76.015 107.78 76.225 108.54 ;
    RECT 76.705 107.78 76.92 108.54 ;
    RECT 77.4 107.78 77.62 108.54 ;
    RECT 78.1 107.78 78.32 108.54 ;
    RECT 78.8 107.78 79.02 108.54 ;
    RECT 79.5 107.78 81.115 108.54 ;
    RECT 81.595 107.78 81.815 108.54 ;
    RECT 82.295 107.78 82.515 108.54 ;
    RECT 82.995 107.78 83.055 108.54 ;
    RECT 83.055 107.69 83.335 108.63 ;
    RECT 83.335 107.78 83.505 108.54 ;
    RECT 26.71 107.02 26.88 107.78 ;
    RECT 26.88 106.93 27.16 107.87 ;
    RECT 27.16 107.02 27.32 107.78 ;
    RECT 27.8 107.02 28.02 107.78 ;
    RECT 28.5 107.02 28.72 107.78 ;
    RECT 29.2 107.02 30.815 107.78 ;
    RECT 31.295 107.02 31.515 107.78 ;
    RECT 31.995 107.02 32.21 107.78 ;
    RECT 32.69 107.02 32.91 107.78 ;
    RECT 33.39 107.02 33.61 107.78 ;
    RECT 34.09 107.02 34.31 107.78 ;
    RECT 34.79 107.02 35.005 107.78 ;
    RECT 35.485 107.02 36.405 107.78 ;
    RECT 36.885 107.02 37.105 107.78 ;
    RECT 37.585 107.02 37.8 107.78 ;
    RECT 38.28 107.02 38.5 107.78 ;
    RECT 38.98 107.02 39.2 107.78 ;
    RECT 39.68 107.02 39.895 107.78 ;
    RECT 40.375 107.02 40.595 107.78 ;
    RECT 41.075 107.02 41.995 107.78 ;
    RECT 42.475 107.02 42.69 107.78 ;
    RECT 43.17 107.02 43.39 107.78 ;
    RECT 43.87 107.02 44.09 107.78 ;
    RECT 44.57 107.02 44.79 107.78 ;
    RECT 45.27 107.02 45.485 107.78 ;
    RECT 45.965 107.02 46.185 107.78 ;
    RECT 46.665 107.02 47.58 107.78 ;
    RECT 48.06 107.02 48.28 107.78 ;
    RECT 48.76 107.02 48.98 107.78 ;
    RECT 49.46 107.02 49.68 107.78 ;
    RECT 50.16 107.02 50.375 107.78 ;
    RECT 50.855 107.02 51.775 107.78 ;
    RECT 52.255 107.02 53.17 107.78 ;
    RECT 53.65 107.02 53.87 107.78 ;
    RECT 54.35 107.02 54.57 107.78 ;
    RECT 55.05 107.02 55.265 107.78 ;
    RECT 55.745 107.02 55.965 107.78 ;
    RECT 56.445 107.02 56.665 107.78 ;
    RECT 57.145 107.02 58.06 107.78 ;
    RECT 58.54 107.02 59.46 107.78 ;
    RECT 59.94 107.02 60.16 107.78 ;
    RECT 60.64 107.02 60.855 107.78 ;
    RECT 61.335 107.02 61.555 107.78 ;
    RECT 62.035 107.02 62.25 107.78 ;
    RECT 62.73 107.02 63.65 107.78 ;
    RECT 64.13 107.02 64.345 107.78 ;
    RECT 64.825 107.02 65.045 107.78 ;
    RECT 65.525 107.02 65.745 107.78 ;
    RECT 66.225 107.02 66.445 107.78 ;
    RECT 66.925 107.02 67.14 107.78 ;
    RECT 67.62 107.02 67.84 107.78 ;
    RECT 68.32 107.02 69.235 107.78 ;
    RECT 69.715 107.02 69.935 107.78 ;
    RECT 70.415 107.02 70.635 107.78 ;
    RECT 71.115 107.02 71.335 107.78 ;
    RECT 71.815 107.02 72.035 107.78 ;
    RECT 72.515 107.02 72.735 107.78 ;
    RECT 73.215 107.02 73.435 107.78 ;
    RECT 73.915 107.02 74.835 107.78 ;
    RECT 75.315 107.02 75.535 107.78 ;
    RECT 76.015 107.02 76.225 107.78 ;
    RECT 76.705 107.02 76.92 107.78 ;
    RECT 77.4 107.02 77.62 107.78 ;
    RECT 78.1 107.02 78.32 107.78 ;
    RECT 78.8 107.02 79.02 107.78 ;
    RECT 79.5 107.02 81.115 107.78 ;
    RECT 81.595 107.02 81.815 107.78 ;
    RECT 82.295 107.02 82.515 107.78 ;
    RECT 82.995 107.02 83.055 107.78 ;
    RECT 83.055 106.93 83.335 107.87 ;
    RECT 83.335 107.02 83.505 107.78 ;
    RECT 26.71 106.26 26.88 107.02 ;
    RECT 26.88 106.17 27.16 107.11 ;
    RECT 27.16 106.26 27.32 107.02 ;
    RECT 27.8 106.26 28.02 107.02 ;
    RECT 28.5 106.26 28.72 107.02 ;
    RECT 29.2 106.26 30.815 107.02 ;
    RECT 31.295 106.26 31.515 107.02 ;
    RECT 31.995 106.26 32.21 107.02 ;
    RECT 32.69 106.26 32.91 107.02 ;
    RECT 33.39 106.26 33.61 107.02 ;
    RECT 34.09 106.26 34.31 107.02 ;
    RECT 34.79 106.26 35.005 107.02 ;
    RECT 35.485 106.26 36.405 107.02 ;
    RECT 36.885 106.26 37.105 107.02 ;
    RECT 37.585 106.26 37.8 107.02 ;
    RECT 38.28 106.26 38.5 107.02 ;
    RECT 38.98 106.26 39.2 107.02 ;
    RECT 39.68 106.26 39.895 107.02 ;
    RECT 40.375 106.26 40.595 107.02 ;
    RECT 41.075 106.26 41.995 107.02 ;
    RECT 42.475 106.26 42.69 107.02 ;
    RECT 43.17 106.26 43.39 107.02 ;
    RECT 43.87 106.26 44.09 107.02 ;
    RECT 44.57 106.26 44.79 107.02 ;
    RECT 45.27 106.26 45.485 107.02 ;
    RECT 45.965 106.26 46.185 107.02 ;
    RECT 46.665 106.26 47.58 107.02 ;
    RECT 48.06 106.26 48.28 107.02 ;
    RECT 48.76 106.26 48.98 107.02 ;
    RECT 49.46 106.26 49.68 107.02 ;
    RECT 50.16 106.26 50.375 107.02 ;
    RECT 50.855 106.26 51.775 107.02 ;
    RECT 52.255 106.26 53.17 107.02 ;
    RECT 53.65 106.26 53.87 107.02 ;
    RECT 54.35 106.26 54.57 107.02 ;
    RECT 55.05 106.26 55.265 107.02 ;
    RECT 55.745 106.26 55.965 107.02 ;
    RECT 56.445 106.26 56.665 107.02 ;
    RECT 57.145 106.26 58.06 107.02 ;
    RECT 58.54 106.26 59.46 107.02 ;
    RECT 59.94 106.26 60.16 107.02 ;
    RECT 60.64 106.26 60.855 107.02 ;
    RECT 61.335 106.26 61.555 107.02 ;
    RECT 62.035 106.26 62.25 107.02 ;
    RECT 62.73 106.26 63.65 107.02 ;
    RECT 64.13 106.26 64.345 107.02 ;
    RECT 64.825 106.26 65.045 107.02 ;
    RECT 65.525 106.26 65.745 107.02 ;
    RECT 66.225 106.26 66.445 107.02 ;
    RECT 66.925 106.26 67.14 107.02 ;
    RECT 67.62 106.26 67.84 107.02 ;
    RECT 68.32 106.26 69.235 107.02 ;
    RECT 69.715 106.26 69.935 107.02 ;
    RECT 70.415 106.26 70.635 107.02 ;
    RECT 71.115 106.26 71.335 107.02 ;
    RECT 71.815 106.26 72.035 107.02 ;
    RECT 72.515 106.26 72.735 107.02 ;
    RECT 73.215 106.26 73.435 107.02 ;
    RECT 73.915 106.26 74.835 107.02 ;
    RECT 75.315 106.26 75.535 107.02 ;
    RECT 76.015 106.26 76.225 107.02 ;
    RECT 76.705 106.26 76.92 107.02 ;
    RECT 77.4 106.26 77.62 107.02 ;
    RECT 78.1 106.26 78.32 107.02 ;
    RECT 78.8 106.26 79.02 107.02 ;
    RECT 79.5 106.26 81.115 107.02 ;
    RECT 81.595 106.26 81.815 107.02 ;
    RECT 82.295 106.26 82.515 107.02 ;
    RECT 82.995 106.26 83.055 107.02 ;
    RECT 83.055 106.17 83.335 107.11 ;
    RECT 83.335 106.26 83.505 107.02 ;
    RECT 26.71 105.5 26.88 106.26 ;
    RECT 26.88 105.41 27.16 106.35 ;
    RECT 27.16 105.5 27.32 106.26 ;
    RECT 27.8 105.5 28.02 106.26 ;
    RECT 28.5 105.5 28.72 106.26 ;
    RECT 29.2 105.5 30.815 106.26 ;
    RECT 31.295 105.5 31.515 106.26 ;
    RECT 31.995 105.5 32.21 106.26 ;
    RECT 32.69 105.5 32.91 106.26 ;
    RECT 33.39 105.5 33.61 106.26 ;
    RECT 34.09 105.5 34.31 106.26 ;
    RECT 34.79 105.5 35.005 106.26 ;
    RECT 35.485 105.5 36.405 106.26 ;
    RECT 36.885 105.5 37.105 106.26 ;
    RECT 37.585 105.5 37.8 106.26 ;
    RECT 38.28 105.5 38.5 106.26 ;
    RECT 38.98 105.5 39.2 106.26 ;
    RECT 39.68 105.5 39.895 106.26 ;
    RECT 40.375 105.5 40.595 106.26 ;
    RECT 41.075 105.5 41.995 106.26 ;
    RECT 42.475 105.5 42.69 106.26 ;
    RECT 43.17 105.5 43.39 106.26 ;
    RECT 43.87 105.5 44.09 106.26 ;
    RECT 44.57 105.5 44.79 106.26 ;
    RECT 45.27 105.5 45.485 106.26 ;
    RECT 45.965 105.5 46.185 106.26 ;
    RECT 46.665 105.5 47.58 106.26 ;
    RECT 48.06 105.5 48.28 106.26 ;
    RECT 48.76 105.5 48.98 106.26 ;
    RECT 49.46 105.5 49.68 106.26 ;
    RECT 50.16 105.5 50.375 106.26 ;
    RECT 50.855 105.5 51.775 106.26 ;
    RECT 52.255 105.5 53.17 106.26 ;
    RECT 53.65 105.5 53.87 106.26 ;
    RECT 54.35 105.5 54.57 106.26 ;
    RECT 55.05 105.5 55.265 106.26 ;
    RECT 55.745 105.5 55.965 106.26 ;
    RECT 56.445 105.5 56.665 106.26 ;
    RECT 57.145 105.5 58.06 106.26 ;
    RECT 58.54 105.5 59.46 106.26 ;
    RECT 59.94 105.5 60.16 106.26 ;
    RECT 60.64 105.5 60.855 106.26 ;
    RECT 61.335 105.5 61.555 106.26 ;
    RECT 62.035 105.5 62.25 106.26 ;
    RECT 62.73 105.5 63.65 106.26 ;
    RECT 64.13 105.5 64.345 106.26 ;
    RECT 64.825 105.5 65.045 106.26 ;
    RECT 65.525 105.5 65.745 106.26 ;
    RECT 66.225 105.5 66.445 106.26 ;
    RECT 66.925 105.5 67.14 106.26 ;
    RECT 67.62 105.5 67.84 106.26 ;
    RECT 68.32 105.5 69.235 106.26 ;
    RECT 69.715 105.5 69.935 106.26 ;
    RECT 70.415 105.5 70.635 106.26 ;
    RECT 71.115 105.5 71.335 106.26 ;
    RECT 71.815 105.5 72.035 106.26 ;
    RECT 72.515 105.5 72.735 106.26 ;
    RECT 73.215 105.5 73.435 106.26 ;
    RECT 73.915 105.5 74.835 106.26 ;
    RECT 75.315 105.5 75.535 106.26 ;
    RECT 76.015 105.5 76.225 106.26 ;
    RECT 76.705 105.5 76.92 106.26 ;
    RECT 77.4 105.5 77.62 106.26 ;
    RECT 78.1 105.5 78.32 106.26 ;
    RECT 78.8 105.5 79.02 106.26 ;
    RECT 79.5 105.5 81.115 106.26 ;
    RECT 81.595 105.5 81.815 106.26 ;
    RECT 82.295 105.5 82.515 106.26 ;
    RECT 82.995 105.5 83.055 106.26 ;
    RECT 83.055 105.41 83.335 106.35 ;
    RECT 83.335 105.5 83.505 106.26 ;
    RECT 26.71 104.74 26.88 105.5 ;
    RECT 26.88 104.65 27.16 105.59 ;
    RECT 27.16 104.74 27.32 105.5 ;
    RECT 27.8 104.74 28.02 105.5 ;
    RECT 28.5 104.74 28.72 105.5 ;
    RECT 29.2 104.74 30.815 105.5 ;
    RECT 31.295 104.74 31.515 105.5 ;
    RECT 31.995 104.74 32.21 105.5 ;
    RECT 32.69 104.74 32.91 105.5 ;
    RECT 33.39 104.74 33.61 105.5 ;
    RECT 34.09 104.74 34.31 105.5 ;
    RECT 34.79 104.74 35.005 105.5 ;
    RECT 35.485 104.74 36.405 105.5 ;
    RECT 36.885 104.74 37.105 105.5 ;
    RECT 37.585 104.74 37.8 105.5 ;
    RECT 38.28 104.74 38.5 105.5 ;
    RECT 38.98 104.74 39.2 105.5 ;
    RECT 39.68 104.74 39.895 105.5 ;
    RECT 40.375 104.74 40.595 105.5 ;
    RECT 41.075 104.74 41.995 105.5 ;
    RECT 42.475 104.74 42.69 105.5 ;
    RECT 43.17 104.74 43.39 105.5 ;
    RECT 43.87 104.74 44.09 105.5 ;
    RECT 44.57 104.74 44.79 105.5 ;
    RECT 45.27 104.74 45.485 105.5 ;
    RECT 45.965 104.74 46.185 105.5 ;
    RECT 46.665 104.74 47.58 105.5 ;
    RECT 48.06 104.74 48.28 105.5 ;
    RECT 48.76 104.74 48.98 105.5 ;
    RECT 49.46 104.74 49.68 105.5 ;
    RECT 50.16 104.74 50.375 105.5 ;
    RECT 50.855 104.74 51.775 105.5 ;
    RECT 52.255 104.74 53.17 105.5 ;
    RECT 53.65 104.74 53.87 105.5 ;
    RECT 54.35 104.74 54.57 105.5 ;
    RECT 55.05 104.74 55.265 105.5 ;
    RECT 55.745 104.74 55.965 105.5 ;
    RECT 56.445 104.74 56.665 105.5 ;
    RECT 57.145 104.74 58.06 105.5 ;
    RECT 58.54 104.74 59.46 105.5 ;
    RECT 59.94 104.74 60.16 105.5 ;
    RECT 60.64 104.74 60.855 105.5 ;
    RECT 61.335 104.74 61.555 105.5 ;
    RECT 62.035 104.74 62.25 105.5 ;
    RECT 62.73 104.74 63.65 105.5 ;
    RECT 64.13 104.74 64.345 105.5 ;
    RECT 64.825 104.74 65.045 105.5 ;
    RECT 65.525 104.74 65.745 105.5 ;
    RECT 66.225 104.74 66.445 105.5 ;
    RECT 66.925 104.74 67.14 105.5 ;
    RECT 67.62 104.74 67.84 105.5 ;
    RECT 68.32 104.74 69.235 105.5 ;
    RECT 69.715 104.74 69.935 105.5 ;
    RECT 70.415 104.74 70.635 105.5 ;
    RECT 71.115 104.74 71.335 105.5 ;
    RECT 71.815 104.74 72.035 105.5 ;
    RECT 72.515 104.74 72.735 105.5 ;
    RECT 73.215 104.74 73.435 105.5 ;
    RECT 73.915 104.74 74.835 105.5 ;
    RECT 75.315 104.74 75.535 105.5 ;
    RECT 76.015 104.74 76.225 105.5 ;
    RECT 76.705 104.74 76.92 105.5 ;
    RECT 77.4 104.74 77.62 105.5 ;
    RECT 78.1 104.74 78.32 105.5 ;
    RECT 78.8 104.74 79.02 105.5 ;
    RECT 79.5 104.74 81.115 105.5 ;
    RECT 81.595 104.74 81.815 105.5 ;
    RECT 82.295 104.74 82.515 105.5 ;
    RECT 82.995 104.74 83.055 105.5 ;
    RECT 83.055 104.65 83.335 105.59 ;
    RECT 83.335 104.74 83.505 105.5 ;
    RECT 26.71 103.98 26.88 104.74 ;
    RECT 26.88 103.89 27.16 104.83 ;
    RECT 27.16 103.98 27.32 104.74 ;
    RECT 27.8 103.98 28.02 104.74 ;
    RECT 28.5 103.98 28.72 104.74 ;
    RECT 29.2 103.98 30.815 104.74 ;
    RECT 31.295 103.98 31.515 104.74 ;
    RECT 31.995 103.98 32.21 104.74 ;
    RECT 32.69 103.98 32.91 104.74 ;
    RECT 33.39 103.98 33.61 104.74 ;
    RECT 34.09 103.98 34.31 104.74 ;
    RECT 34.79 103.98 35.005 104.74 ;
    RECT 35.485 103.98 36.405 104.74 ;
    RECT 36.885 103.98 37.105 104.74 ;
    RECT 37.585 103.98 37.8 104.74 ;
    RECT 38.28 103.98 38.5 104.74 ;
    RECT 38.98 103.98 39.2 104.74 ;
    RECT 39.68 103.98 39.895 104.74 ;
    RECT 40.375 103.98 40.595 104.74 ;
    RECT 41.075 103.98 41.995 104.74 ;
    RECT 42.475 103.98 42.69 104.74 ;
    RECT 43.17 103.98 43.39 104.74 ;
    RECT 43.87 103.98 44.09 104.74 ;
    RECT 44.57 103.98 44.79 104.74 ;
    RECT 45.27 103.98 45.485 104.74 ;
    RECT 45.965 103.98 46.185 104.74 ;
    RECT 46.665 103.98 47.58 104.74 ;
    RECT 48.06 103.98 48.28 104.74 ;
    RECT 48.76 103.98 48.98 104.74 ;
    RECT 49.46 103.98 49.68 104.74 ;
    RECT 50.16 103.98 50.375 104.74 ;
    RECT 50.855 103.98 51.775 104.74 ;
    RECT 52.255 103.98 53.17 104.74 ;
    RECT 53.65 103.98 53.87 104.74 ;
    RECT 54.35 103.98 54.57 104.74 ;
    RECT 55.05 103.98 55.265 104.74 ;
    RECT 55.745 103.98 55.965 104.74 ;
    RECT 56.445 103.98 56.665 104.74 ;
    RECT 57.145 103.98 58.06 104.74 ;
    RECT 58.54 103.98 59.46 104.74 ;
    RECT 59.94 103.98 60.16 104.74 ;
    RECT 60.64 103.98 60.855 104.74 ;
    RECT 61.335 103.98 61.555 104.74 ;
    RECT 62.035 103.98 62.25 104.74 ;
    RECT 62.73 103.98 63.65 104.74 ;
    RECT 64.13 103.98 64.345 104.74 ;
    RECT 64.825 103.98 65.045 104.74 ;
    RECT 65.525 103.98 65.745 104.74 ;
    RECT 66.225 103.98 66.445 104.74 ;
    RECT 66.925 103.98 67.14 104.74 ;
    RECT 67.62 103.98 67.84 104.74 ;
    RECT 68.32 103.98 69.235 104.74 ;
    RECT 69.715 103.98 69.935 104.74 ;
    RECT 70.415 103.98 70.635 104.74 ;
    RECT 71.115 103.98 71.335 104.74 ;
    RECT 71.815 103.98 72.035 104.74 ;
    RECT 72.515 103.98 72.735 104.74 ;
    RECT 73.215 103.98 73.435 104.74 ;
    RECT 73.915 103.98 74.835 104.74 ;
    RECT 75.315 103.98 75.535 104.74 ;
    RECT 76.015 103.98 76.225 104.74 ;
    RECT 76.705 103.98 76.92 104.74 ;
    RECT 77.4 103.98 77.62 104.74 ;
    RECT 78.1 103.98 78.32 104.74 ;
    RECT 78.8 103.98 79.02 104.74 ;
    RECT 79.5 103.98 81.115 104.74 ;
    RECT 81.595 103.98 81.815 104.74 ;
    RECT 82.295 103.98 82.515 104.74 ;
    RECT 82.995 103.98 83.055 104.74 ;
    RECT 83.055 103.89 83.335 104.83 ;
    RECT 83.335 103.98 83.505 104.74 ;
    RECT 26.71 103.22 26.88 103.98 ;
    RECT 26.88 103.13 27.16 104.07 ;
    RECT 27.16 103.22 27.32 103.98 ;
    RECT 27.8 103.22 28.02 103.98 ;
    RECT 28.5 103.22 28.72 103.98 ;
    RECT 29.2 103.22 30.815 103.98 ;
    RECT 31.295 103.22 31.515 103.98 ;
    RECT 31.995 103.22 32.21 103.98 ;
    RECT 32.69 103.22 32.91 103.98 ;
    RECT 33.39 103.22 33.61 103.98 ;
    RECT 34.09 103.22 34.31 103.98 ;
    RECT 34.79 103.22 35.005 103.98 ;
    RECT 35.485 103.22 36.405 103.98 ;
    RECT 36.885 103.22 37.105 103.98 ;
    RECT 37.585 103.22 37.8 103.98 ;
    RECT 38.28 103.22 38.5 103.98 ;
    RECT 38.98 103.22 39.2 103.98 ;
    RECT 39.68 103.22 39.895 103.98 ;
    RECT 40.375 103.22 40.595 103.98 ;
    RECT 41.075 103.22 41.995 103.98 ;
    RECT 42.475 103.22 42.69 103.98 ;
    RECT 43.17 103.22 43.39 103.98 ;
    RECT 43.87 103.22 44.09 103.98 ;
    RECT 44.57 103.22 44.79 103.98 ;
    RECT 45.27 103.22 45.485 103.98 ;
    RECT 45.965 103.22 46.185 103.98 ;
    RECT 46.665 103.22 47.58 103.98 ;
    RECT 48.06 103.22 48.28 103.98 ;
    RECT 48.76 103.22 48.98 103.98 ;
    RECT 49.46 103.22 49.68 103.98 ;
    RECT 50.16 103.22 50.375 103.98 ;
    RECT 50.855 103.22 51.775 103.98 ;
    RECT 52.255 103.22 53.17 103.98 ;
    RECT 53.65 103.22 53.87 103.98 ;
    RECT 54.35 103.22 54.57 103.98 ;
    RECT 55.05 103.22 55.265 103.98 ;
    RECT 55.745 103.22 55.965 103.98 ;
    RECT 56.445 103.22 56.665 103.98 ;
    RECT 57.145 103.22 58.06 103.98 ;
    RECT 58.54 103.22 59.46 103.98 ;
    RECT 59.94 103.22 60.16 103.98 ;
    RECT 60.64 103.22 60.855 103.98 ;
    RECT 61.335 103.22 61.555 103.98 ;
    RECT 62.035 103.22 62.25 103.98 ;
    RECT 62.73 103.22 63.65 103.98 ;
    RECT 64.13 103.22 64.345 103.98 ;
    RECT 64.825 103.22 65.045 103.98 ;
    RECT 65.525 103.22 65.745 103.98 ;
    RECT 66.225 103.22 66.445 103.98 ;
    RECT 66.925 103.22 67.14 103.98 ;
    RECT 67.62 103.22 67.84 103.98 ;
    RECT 68.32 103.22 69.235 103.98 ;
    RECT 69.715 103.22 69.935 103.98 ;
    RECT 70.415 103.22 70.635 103.98 ;
    RECT 71.115 103.22 71.335 103.98 ;
    RECT 71.815 103.22 72.035 103.98 ;
    RECT 72.515 103.22 72.735 103.98 ;
    RECT 73.215 103.22 73.435 103.98 ;
    RECT 73.915 103.22 74.835 103.98 ;
    RECT 75.315 103.22 75.535 103.98 ;
    RECT 76.015 103.22 76.225 103.98 ;
    RECT 76.705 103.22 76.92 103.98 ;
    RECT 77.4 103.22 77.62 103.98 ;
    RECT 78.1 103.22 78.32 103.98 ;
    RECT 78.8 103.22 79.02 103.98 ;
    RECT 79.5 103.22 81.115 103.98 ;
    RECT 81.595 103.22 81.815 103.98 ;
    RECT 82.295 103.22 82.515 103.98 ;
    RECT 82.995 103.22 83.055 103.98 ;
    RECT 83.055 103.13 83.335 104.07 ;
    RECT 83.335 103.22 83.505 103.98 ;
    RECT 26.71 102.46 26.88 103.22 ;
    RECT 26.88 102.37 27.16 103.31 ;
    RECT 27.16 102.46 27.32 103.22 ;
    RECT 27.8 102.46 28.02 103.22 ;
    RECT 28.5 102.46 28.72 103.22 ;
    RECT 29.2 102.46 30.815 103.22 ;
    RECT 31.295 102.46 31.515 103.22 ;
    RECT 31.995 102.46 32.21 103.22 ;
    RECT 32.69 102.46 32.91 103.22 ;
    RECT 33.39 102.46 33.61 103.22 ;
    RECT 34.09 102.46 34.31 103.22 ;
    RECT 34.79 102.46 35.005 103.22 ;
    RECT 35.485 102.46 36.405 103.22 ;
    RECT 36.885 102.46 37.105 103.22 ;
    RECT 37.585 102.46 37.8 103.22 ;
    RECT 38.28 102.46 38.5 103.22 ;
    RECT 38.98 102.46 39.2 103.22 ;
    RECT 39.68 102.46 39.895 103.22 ;
    RECT 40.375 102.46 40.595 103.22 ;
    RECT 41.075 102.46 41.995 103.22 ;
    RECT 42.475 102.46 42.69 103.22 ;
    RECT 43.17 102.46 43.39 103.22 ;
    RECT 43.87 102.46 44.09 103.22 ;
    RECT 44.57 102.46 44.79 103.22 ;
    RECT 45.27 102.46 45.485 103.22 ;
    RECT 45.965 102.46 46.185 103.22 ;
    RECT 46.665 102.46 47.58 103.22 ;
    RECT 48.06 102.46 48.28 103.22 ;
    RECT 48.76 102.46 48.98 103.22 ;
    RECT 49.46 102.46 49.68 103.22 ;
    RECT 50.16 102.46 50.375 103.22 ;
    RECT 50.855 102.46 51.775 103.22 ;
    RECT 52.255 102.46 53.17 103.22 ;
    RECT 53.65 102.46 53.87 103.22 ;
    RECT 54.35 102.46 54.57 103.22 ;
    RECT 55.05 102.46 55.265 103.22 ;
    RECT 55.745 102.46 55.965 103.22 ;
    RECT 56.445 102.46 56.665 103.22 ;
    RECT 57.145 102.46 58.06 103.22 ;
    RECT 58.54 102.46 59.46 103.22 ;
    RECT 59.94 102.46 60.16 103.22 ;
    RECT 60.64 102.46 60.855 103.22 ;
    RECT 61.335 102.46 61.555 103.22 ;
    RECT 62.035 102.46 62.25 103.22 ;
    RECT 62.73 102.46 63.65 103.22 ;
    RECT 64.13 102.46 64.345 103.22 ;
    RECT 64.825 102.46 65.045 103.22 ;
    RECT 65.525 102.46 65.745 103.22 ;
    RECT 66.225 102.46 66.445 103.22 ;
    RECT 66.925 102.46 67.14 103.22 ;
    RECT 67.62 102.46 67.84 103.22 ;
    RECT 68.32 102.46 69.235 103.22 ;
    RECT 69.715 102.46 69.935 103.22 ;
    RECT 70.415 102.46 70.635 103.22 ;
    RECT 71.115 102.46 71.335 103.22 ;
    RECT 71.815 102.46 72.035 103.22 ;
    RECT 72.515 102.46 72.735 103.22 ;
    RECT 73.215 102.46 73.435 103.22 ;
    RECT 73.915 102.46 74.835 103.22 ;
    RECT 75.315 102.46 75.535 103.22 ;
    RECT 76.015 102.46 76.225 103.22 ;
    RECT 76.705 102.46 76.92 103.22 ;
    RECT 77.4 102.46 77.62 103.22 ;
    RECT 78.1 102.46 78.32 103.22 ;
    RECT 78.8 102.46 79.02 103.22 ;
    RECT 79.5 102.46 81.115 103.22 ;
    RECT 81.595 102.46 81.815 103.22 ;
    RECT 82.295 102.46 82.515 103.22 ;
    RECT 82.995 102.46 83.055 103.22 ;
    RECT 83.055 102.37 83.335 103.31 ;
    RECT 83.335 102.46 83.505 103.22 ;
    RECT 26.71 101.7 26.88 102.46 ;
    RECT 26.88 101.61 27.16 102.55 ;
    RECT 27.16 101.7 27.32 102.46 ;
    RECT 27.8 101.7 28.02 102.46 ;
    RECT 28.5 101.7 28.72 102.46 ;
    RECT 29.2 101.7 30.815 102.46 ;
    RECT 31.295 101.7 31.515 102.46 ;
    RECT 31.995 101.7 32.21 102.46 ;
    RECT 32.69 101.7 32.91 102.46 ;
    RECT 33.39 101.7 33.61 102.46 ;
    RECT 34.09 101.7 34.31 102.46 ;
    RECT 34.79 101.7 35.005 102.46 ;
    RECT 35.485 101.7 36.405 102.46 ;
    RECT 36.885 101.7 37.105 102.46 ;
    RECT 37.585 101.7 37.8 102.46 ;
    RECT 38.28 101.7 38.5 102.46 ;
    RECT 38.98 101.7 39.2 102.46 ;
    RECT 39.68 101.7 39.895 102.46 ;
    RECT 40.375 101.7 40.595 102.46 ;
    RECT 41.075 101.7 41.995 102.46 ;
    RECT 42.475 101.7 42.69 102.46 ;
    RECT 43.17 101.7 43.39 102.46 ;
    RECT 43.87 101.7 44.09 102.46 ;
    RECT 44.57 101.7 44.79 102.46 ;
    RECT 45.27 101.7 45.485 102.46 ;
    RECT 45.965 101.7 46.185 102.46 ;
    RECT 46.665 101.7 47.58 102.46 ;
    RECT 48.06 101.7 48.28 102.46 ;
    RECT 48.76 101.7 48.98 102.46 ;
    RECT 49.46 101.7 49.68 102.46 ;
    RECT 50.16 101.7 50.375 102.46 ;
    RECT 50.855 101.7 51.775 102.46 ;
    RECT 52.255 101.7 53.17 102.46 ;
    RECT 53.65 101.7 53.87 102.46 ;
    RECT 54.35 101.7 54.57 102.46 ;
    RECT 55.05 101.7 55.265 102.46 ;
    RECT 55.745 101.7 55.965 102.46 ;
    RECT 56.445 101.7 56.665 102.46 ;
    RECT 57.145 101.7 58.06 102.46 ;
    RECT 58.54 101.7 59.46 102.46 ;
    RECT 59.94 101.7 60.16 102.46 ;
    RECT 60.64 101.7 60.855 102.46 ;
    RECT 61.335 101.7 61.555 102.46 ;
    RECT 62.035 101.7 62.25 102.46 ;
    RECT 62.73 101.7 63.65 102.46 ;
    RECT 64.13 101.7 64.345 102.46 ;
    RECT 64.825 101.7 65.045 102.46 ;
    RECT 65.525 101.7 65.745 102.46 ;
    RECT 66.225 101.7 66.445 102.46 ;
    RECT 66.925 101.7 67.14 102.46 ;
    RECT 67.62 101.7 67.84 102.46 ;
    RECT 68.32 101.7 69.235 102.46 ;
    RECT 69.715 101.7 69.935 102.46 ;
    RECT 70.415 101.7 70.635 102.46 ;
    RECT 71.115 101.7 71.335 102.46 ;
    RECT 71.815 101.7 72.035 102.46 ;
    RECT 72.515 101.7 72.735 102.46 ;
    RECT 73.215 101.7 73.435 102.46 ;
    RECT 73.915 101.7 74.835 102.46 ;
    RECT 75.315 101.7 75.535 102.46 ;
    RECT 76.015 101.7 76.225 102.46 ;
    RECT 76.705 101.7 76.92 102.46 ;
    RECT 77.4 101.7 77.62 102.46 ;
    RECT 78.1 101.7 78.32 102.46 ;
    RECT 78.8 101.7 79.02 102.46 ;
    RECT 79.5 101.7 81.115 102.46 ;
    RECT 81.595 101.7 81.815 102.46 ;
    RECT 82.295 101.7 82.515 102.46 ;
    RECT 82.995 101.7 83.055 102.46 ;
    RECT 83.055 101.61 83.335 102.55 ;
    RECT 83.335 101.7 83.505 102.46 ;
    RECT 26.71 100.94 26.88 101.7 ;
    RECT 26.88 100.85 27.16 101.79 ;
    RECT 27.16 100.94 27.32 101.7 ;
    RECT 27.8 100.94 28.02 101.7 ;
    RECT 28.5 100.94 28.72 101.7 ;
    RECT 29.2 100.94 30.815 101.7 ;
    RECT 31.295 100.94 31.515 101.7 ;
    RECT 31.995 100.94 32.21 101.7 ;
    RECT 32.69 100.94 32.91 101.7 ;
    RECT 33.39 100.94 33.61 101.7 ;
    RECT 34.09 100.94 34.31 101.7 ;
    RECT 34.79 100.94 35.005 101.7 ;
    RECT 35.485 100.94 36.405 101.7 ;
    RECT 36.885 100.94 37.105 101.7 ;
    RECT 37.585 100.94 37.8 101.7 ;
    RECT 38.28 100.94 38.5 101.7 ;
    RECT 38.98 100.94 39.2 101.7 ;
    RECT 39.68 100.94 39.895 101.7 ;
    RECT 40.375 100.94 40.595 101.7 ;
    RECT 41.075 100.94 41.995 101.7 ;
    RECT 42.475 100.94 42.69 101.7 ;
    RECT 43.17 100.94 43.39 101.7 ;
    RECT 43.87 100.94 44.09 101.7 ;
    RECT 44.57 100.94 44.79 101.7 ;
    RECT 45.27 100.94 45.485 101.7 ;
    RECT 45.965 100.94 46.185 101.7 ;
    RECT 46.665 100.94 47.58 101.7 ;
    RECT 48.06 100.94 48.28 101.7 ;
    RECT 48.76 100.94 48.98 101.7 ;
    RECT 49.46 100.94 49.68 101.7 ;
    RECT 50.16 100.94 50.375 101.7 ;
    RECT 50.855 100.94 51.775 101.7 ;
    RECT 52.255 100.94 53.17 101.7 ;
    RECT 53.65 100.94 53.87 101.7 ;
    RECT 54.35 100.94 54.57 101.7 ;
    RECT 55.05 100.94 55.265 101.7 ;
    RECT 55.745 100.94 55.965 101.7 ;
    RECT 56.445 100.94 56.665 101.7 ;
    RECT 57.145 100.94 58.06 101.7 ;
    RECT 58.54 100.94 59.46 101.7 ;
    RECT 59.94 100.94 60.16 101.7 ;
    RECT 60.64 100.94 60.855 101.7 ;
    RECT 61.335 100.94 61.555 101.7 ;
    RECT 62.035 100.94 62.25 101.7 ;
    RECT 62.73 100.94 63.65 101.7 ;
    RECT 64.13 100.94 64.345 101.7 ;
    RECT 64.825 100.94 65.045 101.7 ;
    RECT 65.525 100.94 65.745 101.7 ;
    RECT 66.225 100.94 66.445 101.7 ;
    RECT 66.925 100.94 67.14 101.7 ;
    RECT 67.62 100.94 67.84 101.7 ;
    RECT 68.32 100.94 69.235 101.7 ;
    RECT 69.715 100.94 69.935 101.7 ;
    RECT 70.415 100.94 70.635 101.7 ;
    RECT 71.115 100.94 71.335 101.7 ;
    RECT 71.815 100.94 72.035 101.7 ;
    RECT 72.515 100.94 72.735 101.7 ;
    RECT 73.215 100.94 73.435 101.7 ;
    RECT 73.915 100.94 74.835 101.7 ;
    RECT 75.315 100.94 75.535 101.7 ;
    RECT 76.015 100.94 76.225 101.7 ;
    RECT 76.705 100.94 76.92 101.7 ;
    RECT 77.4 100.94 77.62 101.7 ;
    RECT 78.1 100.94 78.32 101.7 ;
    RECT 78.8 100.94 79.02 101.7 ;
    RECT 79.5 100.94 81.115 101.7 ;
    RECT 81.595 100.94 81.815 101.7 ;
    RECT 82.295 100.94 82.515 101.7 ;
    RECT 82.995 100.94 83.055 101.7 ;
    RECT 83.055 100.85 83.335 101.79 ;
    RECT 83.335 100.94 83.505 101.7 ;
    RECT 26.71 100.18 26.88 100.94 ;
    RECT 26.88 100.09 27.16 101.03 ;
    RECT 27.16 100.18 27.32 100.94 ;
    RECT 27.8 100.18 28.02 100.94 ;
    RECT 28.5 100.18 28.72 100.94 ;
    RECT 29.2 100.18 30.815 100.94 ;
    RECT 31.295 100.18 31.515 100.94 ;
    RECT 31.995 100.18 32.21 100.94 ;
    RECT 32.69 100.18 32.91 100.94 ;
    RECT 33.39 100.18 33.61 100.94 ;
    RECT 34.09 100.18 34.31 100.94 ;
    RECT 34.79 100.18 35.005 100.94 ;
    RECT 35.485 100.18 36.405 100.94 ;
    RECT 36.885 100.18 37.105 100.94 ;
    RECT 37.585 100.18 37.8 100.94 ;
    RECT 38.28 100.18 38.5 100.94 ;
    RECT 38.98 100.18 39.2 100.94 ;
    RECT 39.68 100.18 39.895 100.94 ;
    RECT 40.375 100.18 40.595 100.94 ;
    RECT 41.075 100.18 41.995 100.94 ;
    RECT 42.475 100.18 42.69 100.94 ;
    RECT 43.17 100.18 43.39 100.94 ;
    RECT 43.87 100.18 44.09 100.94 ;
    RECT 44.57 100.18 44.79 100.94 ;
    RECT 45.27 100.18 45.485 100.94 ;
    RECT 45.965 100.18 46.185 100.94 ;
    RECT 46.665 100.18 47.58 100.94 ;
    RECT 48.06 100.18 48.28 100.94 ;
    RECT 48.76 100.18 48.98 100.94 ;
    RECT 49.46 100.18 49.68 100.94 ;
    RECT 50.16 100.18 50.375 100.94 ;
    RECT 50.855 100.18 51.775 100.94 ;
    RECT 52.255 100.18 53.17 100.94 ;
    RECT 53.65 100.18 53.87 100.94 ;
    RECT 54.35 100.18 54.57 100.94 ;
    RECT 55.05 100.18 55.265 100.94 ;
    RECT 55.745 100.18 55.965 100.94 ;
    RECT 56.445 100.18 56.665 100.94 ;
    RECT 57.145 100.18 58.06 100.94 ;
    RECT 58.54 100.18 59.46 100.94 ;
    RECT 59.94 100.18 60.16 100.94 ;
    RECT 60.64 100.18 60.855 100.94 ;
    RECT 61.335 100.18 61.555 100.94 ;
    RECT 62.035 100.18 62.25 100.94 ;
    RECT 62.73 100.18 63.65 100.94 ;
    RECT 64.13 100.18 64.345 100.94 ;
    RECT 64.825 100.18 65.045 100.94 ;
    RECT 65.525 100.18 65.745 100.94 ;
    RECT 66.225 100.18 66.445 100.94 ;
    RECT 66.925 100.18 67.14 100.94 ;
    RECT 67.62 100.18 67.84 100.94 ;
    RECT 68.32 100.18 69.235 100.94 ;
    RECT 69.715 100.18 69.935 100.94 ;
    RECT 70.415 100.18 70.635 100.94 ;
    RECT 71.115 100.18 71.335 100.94 ;
    RECT 71.815 100.18 72.035 100.94 ;
    RECT 72.515 100.18 72.735 100.94 ;
    RECT 73.215 100.18 73.435 100.94 ;
    RECT 73.915 100.18 74.835 100.94 ;
    RECT 75.315 100.18 75.535 100.94 ;
    RECT 76.015 100.18 76.225 100.94 ;
    RECT 76.705 100.18 76.92 100.94 ;
    RECT 77.4 100.18 77.62 100.94 ;
    RECT 78.1 100.18 78.32 100.94 ;
    RECT 78.8 100.18 79.02 100.94 ;
    RECT 79.5 100.18 81.115 100.94 ;
    RECT 81.595 100.18 81.815 100.94 ;
    RECT 82.295 100.18 82.515 100.94 ;
    RECT 82.995 100.18 83.055 100.94 ;
    RECT 83.055 100.09 83.335 101.03 ;
    RECT 83.335 100.18 83.505 100.94 ;
    RECT 26.71 99.42 26.88 100.18 ;
    RECT 26.88 99.33 27.16 100.27 ;
    RECT 27.16 99.42 27.32 100.18 ;
    RECT 27.8 99.42 28.02 100.18 ;
    RECT 28.5 99.42 28.72 100.18 ;
    RECT 29.2 99.42 30.815 100.18 ;
    RECT 31.295 99.42 31.515 100.18 ;
    RECT 31.995 99.42 32.21 100.18 ;
    RECT 32.69 99.42 32.91 100.18 ;
    RECT 33.39 99.42 33.61 100.18 ;
    RECT 34.09 99.42 34.31 100.18 ;
    RECT 34.79 99.42 35.005 100.18 ;
    RECT 35.485 99.42 36.405 100.18 ;
    RECT 36.885 99.42 37.105 100.18 ;
    RECT 37.585 99.42 37.8 100.18 ;
    RECT 38.28 99.42 38.5 100.18 ;
    RECT 38.98 99.42 39.2 100.18 ;
    RECT 39.68 99.42 39.895 100.18 ;
    RECT 40.375 99.42 40.595 100.18 ;
    RECT 41.075 99.42 41.995 100.18 ;
    RECT 42.475 99.42 42.69 100.18 ;
    RECT 43.17 99.42 43.39 100.18 ;
    RECT 43.87 99.42 44.09 100.18 ;
    RECT 44.57 99.42 44.79 100.18 ;
    RECT 45.27 99.42 45.485 100.18 ;
    RECT 45.965 99.42 46.185 100.18 ;
    RECT 46.665 99.42 47.58 100.18 ;
    RECT 48.06 99.42 48.28 100.18 ;
    RECT 48.76 99.42 48.98 100.18 ;
    RECT 49.46 99.42 49.68 100.18 ;
    RECT 50.16 99.42 50.375 100.18 ;
    RECT 50.855 99.42 51.775 100.18 ;
    RECT 52.255 99.42 53.17 100.18 ;
    RECT 53.65 99.42 53.87 100.18 ;
    RECT 54.35 99.42 54.57 100.18 ;
    RECT 55.05 99.42 55.265 100.18 ;
    RECT 55.745 99.42 55.965 100.18 ;
    RECT 56.445 99.42 56.665 100.18 ;
    RECT 57.145 99.42 58.06 100.18 ;
    RECT 58.54 99.42 59.46 100.18 ;
    RECT 59.94 99.42 60.16 100.18 ;
    RECT 60.64 99.42 60.855 100.18 ;
    RECT 61.335 99.42 61.555 100.18 ;
    RECT 62.035 99.42 62.25 100.18 ;
    RECT 62.73 99.42 63.65 100.18 ;
    RECT 64.13 99.42 64.345 100.18 ;
    RECT 64.825 99.42 65.045 100.18 ;
    RECT 65.525 99.42 65.745 100.18 ;
    RECT 66.225 99.42 66.445 100.18 ;
    RECT 66.925 99.42 67.14 100.18 ;
    RECT 67.62 99.42 67.84 100.18 ;
    RECT 68.32 99.42 69.235 100.18 ;
    RECT 69.715 99.42 69.935 100.18 ;
    RECT 70.415 99.42 70.635 100.18 ;
    RECT 71.115 99.42 71.335 100.18 ;
    RECT 71.815 99.42 72.035 100.18 ;
    RECT 72.515 99.42 72.735 100.18 ;
    RECT 73.215 99.42 73.435 100.18 ;
    RECT 73.915 99.42 74.835 100.18 ;
    RECT 75.315 99.42 75.535 100.18 ;
    RECT 76.015 99.42 76.225 100.18 ;
    RECT 76.705 99.42 76.92 100.18 ;
    RECT 77.4 99.42 77.62 100.18 ;
    RECT 78.1 99.42 78.32 100.18 ;
    RECT 78.8 99.42 79.02 100.18 ;
    RECT 79.5 99.42 81.115 100.18 ;
    RECT 81.595 99.42 81.815 100.18 ;
    RECT 82.295 99.42 82.515 100.18 ;
    RECT 82.995 99.42 83.055 100.18 ;
    RECT 83.055 99.33 83.335 100.27 ;
    RECT 83.335 99.42 83.505 100.18 ;
    RECT 26.71 98.66 26.88 99.42 ;
    RECT 26.88 98.57 27.16 99.51 ;
    RECT 27.16 98.66 27.32 99.42 ;
    RECT 27.8 98.66 28.02 99.42 ;
    RECT 28.5 98.66 28.72 99.42 ;
    RECT 29.2 98.66 30.815 99.42 ;
    RECT 31.295 98.66 31.515 99.42 ;
    RECT 31.995 98.66 32.21 99.42 ;
    RECT 32.69 98.66 32.91 99.42 ;
    RECT 33.39 98.66 33.61 99.42 ;
    RECT 34.09 98.66 34.31 99.42 ;
    RECT 34.79 98.66 35.005 99.42 ;
    RECT 35.485 98.66 36.405 99.42 ;
    RECT 36.885 98.66 37.105 99.42 ;
    RECT 37.585 98.66 37.8 99.42 ;
    RECT 38.28 98.66 38.5 99.42 ;
    RECT 38.98 98.66 39.2 99.42 ;
    RECT 39.68 98.66 39.895 99.42 ;
    RECT 40.375 98.66 40.595 99.42 ;
    RECT 41.075 98.66 41.995 99.42 ;
    RECT 42.475 98.66 42.69 99.42 ;
    RECT 43.17 98.66 43.39 99.42 ;
    RECT 43.87 98.66 44.09 99.42 ;
    RECT 44.57 98.66 44.79 99.42 ;
    RECT 45.27 98.66 45.485 99.42 ;
    RECT 45.965 98.66 46.185 99.42 ;
    RECT 46.665 98.66 47.58 99.42 ;
    RECT 48.06 98.66 48.28 99.42 ;
    RECT 48.76 98.66 48.98 99.42 ;
    RECT 49.46 98.66 49.68 99.42 ;
    RECT 50.16 98.66 50.375 99.42 ;
    RECT 50.855 98.66 51.775 99.42 ;
    RECT 52.255 98.66 53.17 99.42 ;
    RECT 53.65 98.66 53.87 99.42 ;
    RECT 54.35 98.66 54.57 99.42 ;
    RECT 55.05 98.66 55.265 99.42 ;
    RECT 55.745 98.66 55.965 99.42 ;
    RECT 56.445 98.66 56.665 99.42 ;
    RECT 57.145 98.66 58.06 99.42 ;
    RECT 58.54 98.66 59.46 99.42 ;
    RECT 59.94 98.66 60.16 99.42 ;
    RECT 60.64 98.66 60.855 99.42 ;
    RECT 61.335 98.66 61.555 99.42 ;
    RECT 62.035 98.66 62.25 99.42 ;
    RECT 62.73 98.66 63.65 99.42 ;
    RECT 64.13 98.66 64.345 99.42 ;
    RECT 64.825 98.66 65.045 99.42 ;
    RECT 65.525 98.66 65.745 99.42 ;
    RECT 66.225 98.66 66.445 99.42 ;
    RECT 66.925 98.66 67.14 99.42 ;
    RECT 67.62 98.66 67.84 99.42 ;
    RECT 68.32 98.66 69.235 99.42 ;
    RECT 69.715 98.66 69.935 99.42 ;
    RECT 70.415 98.66 70.635 99.42 ;
    RECT 71.115 98.66 71.335 99.42 ;
    RECT 71.815 98.66 72.035 99.42 ;
    RECT 72.515 98.66 72.735 99.42 ;
    RECT 73.215 98.66 73.435 99.42 ;
    RECT 73.915 98.66 74.835 99.42 ;
    RECT 75.315 98.66 75.535 99.42 ;
    RECT 76.015 98.66 76.225 99.42 ;
    RECT 76.705 98.66 76.92 99.42 ;
    RECT 77.4 98.66 77.62 99.42 ;
    RECT 78.1 98.66 78.32 99.42 ;
    RECT 78.8 98.66 79.02 99.42 ;
    RECT 79.5 98.66 81.115 99.42 ;
    RECT 81.595 98.66 81.815 99.42 ;
    RECT 82.295 98.66 82.515 99.42 ;
    RECT 82.995 98.66 83.055 99.42 ;
    RECT 83.055 98.57 83.335 99.51 ;
    RECT 83.335 98.66 83.505 99.42 ;
    RECT 26.71 97.9 26.88 98.66 ;
    RECT 26.88 97.81 27.16 98.75 ;
    RECT 27.16 97.9 27.32 98.66 ;
    RECT 27.8 97.9 28.02 98.66 ;
    RECT 28.5 97.9 28.72 98.66 ;
    RECT 29.2 97.9 30.815 98.66 ;
    RECT 31.295 97.9 31.515 98.66 ;
    RECT 31.995 97.9 32.21 98.66 ;
    RECT 32.69 97.9 32.91 98.66 ;
    RECT 33.39 97.9 33.61 98.66 ;
    RECT 34.09 97.9 34.31 98.66 ;
    RECT 34.79 97.9 35.005 98.66 ;
    RECT 35.485 97.9 36.405 98.66 ;
    RECT 36.885 97.9 37.105 98.66 ;
    RECT 37.585 97.9 37.8 98.66 ;
    RECT 38.28 97.9 38.5 98.66 ;
    RECT 38.98 97.9 39.2 98.66 ;
    RECT 39.68 97.9 39.895 98.66 ;
    RECT 40.375 97.9 40.595 98.66 ;
    RECT 41.075 97.9 41.995 98.66 ;
    RECT 42.475 97.9 42.69 98.66 ;
    RECT 43.17 97.9 43.39 98.66 ;
    RECT 43.87 97.9 44.09 98.66 ;
    RECT 44.57 97.9 44.79 98.66 ;
    RECT 45.27 97.9 45.485 98.66 ;
    RECT 45.965 97.9 46.185 98.66 ;
    RECT 46.665 97.9 47.58 98.66 ;
    RECT 48.06 97.9 48.28 98.66 ;
    RECT 48.76 97.9 48.98 98.66 ;
    RECT 49.46 97.9 49.68 98.66 ;
    RECT 50.16 97.9 50.375 98.66 ;
    RECT 50.855 97.9 51.775 98.66 ;
    RECT 52.255 97.9 53.17 98.66 ;
    RECT 53.65 97.9 53.87 98.66 ;
    RECT 54.35 97.9 54.57 98.66 ;
    RECT 55.05 97.9 55.265 98.66 ;
    RECT 55.745 97.9 55.965 98.66 ;
    RECT 56.445 97.9 56.665 98.66 ;
    RECT 57.145 97.9 58.06 98.66 ;
    RECT 58.54 97.9 59.46 98.66 ;
    RECT 59.94 97.9 60.16 98.66 ;
    RECT 60.64 97.9 60.855 98.66 ;
    RECT 61.335 97.9 61.555 98.66 ;
    RECT 62.035 97.9 62.25 98.66 ;
    RECT 62.73 97.9 63.65 98.66 ;
    RECT 64.13 97.9 64.345 98.66 ;
    RECT 64.825 97.9 65.045 98.66 ;
    RECT 65.525 97.9 65.745 98.66 ;
    RECT 66.225 97.9 66.445 98.66 ;
    RECT 66.925 97.9 67.14 98.66 ;
    RECT 67.62 97.9 67.84 98.66 ;
    RECT 68.32 97.9 69.235 98.66 ;
    RECT 69.715 97.9 69.935 98.66 ;
    RECT 70.415 97.9 70.635 98.66 ;
    RECT 71.115 97.9 71.335 98.66 ;
    RECT 71.815 97.9 72.035 98.66 ;
    RECT 72.515 97.9 72.735 98.66 ;
    RECT 73.215 97.9 73.435 98.66 ;
    RECT 73.915 97.9 74.835 98.66 ;
    RECT 75.315 97.9 75.535 98.66 ;
    RECT 76.015 97.9 76.225 98.66 ;
    RECT 76.705 97.9 76.92 98.66 ;
    RECT 77.4 97.9 77.62 98.66 ;
    RECT 78.1 97.9 78.32 98.66 ;
    RECT 78.8 97.9 79.02 98.66 ;
    RECT 79.5 97.9 81.115 98.66 ;
    RECT 81.595 97.9 81.815 98.66 ;
    RECT 82.295 97.9 82.515 98.66 ;
    RECT 82.995 97.9 83.055 98.66 ;
    RECT 83.055 97.81 83.335 98.75 ;
    RECT 83.335 97.9 83.505 98.66 ;
    RECT 26.71 97.14 26.88 97.9 ;
    RECT 26.88 97.05 27.16 97.99 ;
    RECT 27.16 97.14 27.32 97.9 ;
    RECT 27.8 97.14 28.02 97.9 ;
    RECT 28.5 97.14 28.72 97.9 ;
    RECT 29.2 97.14 30.815 97.9 ;
    RECT 31.295 97.14 31.515 97.9 ;
    RECT 31.995 97.14 32.21 97.9 ;
    RECT 32.69 97.14 32.91 97.9 ;
    RECT 33.39 97.14 33.61 97.9 ;
    RECT 34.09 97.14 34.31 97.9 ;
    RECT 34.79 97.14 35.005 97.9 ;
    RECT 35.485 97.14 36.405 97.9 ;
    RECT 36.885 97.14 37.105 97.9 ;
    RECT 37.585 97.14 37.8 97.9 ;
    RECT 38.28 97.14 38.5 97.9 ;
    RECT 38.98 97.14 39.2 97.9 ;
    RECT 39.68 97.14 39.895 97.9 ;
    RECT 40.375 97.14 40.595 97.9 ;
    RECT 41.075 97.14 41.995 97.9 ;
    RECT 42.475 97.14 42.69 97.9 ;
    RECT 43.17 97.14 43.39 97.9 ;
    RECT 43.87 97.14 44.09 97.9 ;
    RECT 44.57 97.14 44.79 97.9 ;
    RECT 45.27 97.14 45.485 97.9 ;
    RECT 45.965 97.14 46.185 97.9 ;
    RECT 46.665 97.14 47.58 97.9 ;
    RECT 48.06 97.14 48.28 97.9 ;
    RECT 48.76 97.14 48.98 97.9 ;
    RECT 49.46 97.14 49.68 97.9 ;
    RECT 50.16 97.14 50.375 97.9 ;
    RECT 50.855 97.14 51.775 97.9 ;
    RECT 52.255 97.14 53.17 97.9 ;
    RECT 53.65 97.14 53.87 97.9 ;
    RECT 54.35 97.14 54.57 97.9 ;
    RECT 55.05 97.14 55.265 97.9 ;
    RECT 55.745 97.14 55.965 97.9 ;
    RECT 56.445 97.14 56.665 97.9 ;
    RECT 57.145 97.14 58.06 97.9 ;
    RECT 58.54 97.14 59.46 97.9 ;
    RECT 59.94 97.14 60.16 97.9 ;
    RECT 60.64 97.14 60.855 97.9 ;
    RECT 61.335 97.14 61.555 97.9 ;
    RECT 62.035 97.14 62.25 97.9 ;
    RECT 62.73 97.14 63.65 97.9 ;
    RECT 64.13 97.14 64.345 97.9 ;
    RECT 64.825 97.14 65.045 97.9 ;
    RECT 65.525 97.14 65.745 97.9 ;
    RECT 66.225 97.14 66.445 97.9 ;
    RECT 66.925 97.14 67.14 97.9 ;
    RECT 67.62 97.14 67.84 97.9 ;
    RECT 68.32 97.14 69.235 97.9 ;
    RECT 69.715 97.14 69.935 97.9 ;
    RECT 70.415 97.14 70.635 97.9 ;
    RECT 71.115 97.14 71.335 97.9 ;
    RECT 71.815 97.14 72.035 97.9 ;
    RECT 72.515 97.14 72.735 97.9 ;
    RECT 73.215 97.14 73.435 97.9 ;
    RECT 73.915 97.14 74.835 97.9 ;
    RECT 75.315 97.14 75.535 97.9 ;
    RECT 76.015 97.14 76.225 97.9 ;
    RECT 76.705 97.14 76.92 97.9 ;
    RECT 77.4 97.14 77.62 97.9 ;
    RECT 78.1 97.14 78.32 97.9 ;
    RECT 78.8 97.14 79.02 97.9 ;
    RECT 79.5 97.14 81.115 97.9 ;
    RECT 81.595 97.14 81.815 97.9 ;
    RECT 82.295 97.14 82.515 97.9 ;
    RECT 82.995 97.14 83.055 97.9 ;
    RECT 83.055 97.05 83.335 97.99 ;
    RECT 83.335 97.14 83.505 97.9 ;
    RECT 26.71 96.38 26.88 97.14 ;
    RECT 26.88 96.29 27.16 97.23 ;
    RECT 27.16 96.38 27.32 97.14 ;
    RECT 27.8 96.38 28.02 97.14 ;
    RECT 28.5 96.38 28.72 97.14 ;
    RECT 29.2 96.38 30.815 97.14 ;
    RECT 31.295 96.38 31.515 97.14 ;
    RECT 31.995 96.38 32.21 97.14 ;
    RECT 32.69 96.38 32.91 97.14 ;
    RECT 33.39 96.38 33.61 97.14 ;
    RECT 34.09 96.38 34.31 97.14 ;
    RECT 34.79 96.38 35.005 97.14 ;
    RECT 35.485 96.38 36.405 97.14 ;
    RECT 36.885 96.38 37.105 97.14 ;
    RECT 37.585 96.38 37.8 97.14 ;
    RECT 38.28 96.38 38.5 97.14 ;
    RECT 38.98 96.38 39.2 97.14 ;
    RECT 39.68 96.38 39.895 97.14 ;
    RECT 40.375 96.38 40.595 97.14 ;
    RECT 41.075 96.38 41.995 97.14 ;
    RECT 42.475 96.38 42.69 97.14 ;
    RECT 43.17 96.38 43.39 97.14 ;
    RECT 43.87 96.38 44.09 97.14 ;
    RECT 44.57 96.38 44.79 97.14 ;
    RECT 45.27 96.38 45.485 97.14 ;
    RECT 45.965 96.38 46.185 97.14 ;
    RECT 46.665 96.38 47.58 97.14 ;
    RECT 48.06 96.38 48.28 97.14 ;
    RECT 48.76 96.38 48.98 97.14 ;
    RECT 49.46 96.38 49.68 97.14 ;
    RECT 50.16 96.38 50.375 97.14 ;
    RECT 50.855 96.38 51.775 97.14 ;
    RECT 52.255 96.38 53.17 97.14 ;
    RECT 53.65 96.38 53.87 97.14 ;
    RECT 54.35 96.38 54.57 97.14 ;
    RECT 55.05 96.38 55.265 97.14 ;
    RECT 55.745 96.38 55.965 97.14 ;
    RECT 56.445 96.38 56.665 97.14 ;
    RECT 57.145 96.38 58.06 97.14 ;
    RECT 58.54 96.38 59.46 97.14 ;
    RECT 59.94 96.38 60.16 97.14 ;
    RECT 60.64 96.38 60.855 97.14 ;
    RECT 61.335 96.38 61.555 97.14 ;
    RECT 62.035 96.38 62.25 97.14 ;
    RECT 62.73 96.38 63.65 97.14 ;
    RECT 64.13 96.38 64.345 97.14 ;
    RECT 64.825 96.38 65.045 97.14 ;
    RECT 65.525 96.38 65.745 97.14 ;
    RECT 66.225 96.38 66.445 97.14 ;
    RECT 66.925 96.38 67.14 97.14 ;
    RECT 67.62 96.38 67.84 97.14 ;
    RECT 68.32 96.38 69.235 97.14 ;
    RECT 69.715 96.38 69.935 97.14 ;
    RECT 70.415 96.38 70.635 97.14 ;
    RECT 71.115 96.38 71.335 97.14 ;
    RECT 71.815 96.38 72.035 97.14 ;
    RECT 72.515 96.38 72.735 97.14 ;
    RECT 73.215 96.38 73.435 97.14 ;
    RECT 73.915 96.38 74.835 97.14 ;
    RECT 75.315 96.38 75.535 97.14 ;
    RECT 76.015 96.38 76.225 97.14 ;
    RECT 76.705 96.38 76.92 97.14 ;
    RECT 77.4 96.38 77.62 97.14 ;
    RECT 78.1 96.38 78.32 97.14 ;
    RECT 78.8 96.38 79.02 97.14 ;
    RECT 79.5 96.38 81.115 97.14 ;
    RECT 81.595 96.38 81.815 97.14 ;
    RECT 82.295 96.38 82.515 97.14 ;
    RECT 82.995 96.38 83.055 97.14 ;
    RECT 83.055 96.29 83.335 97.23 ;
    RECT 83.335 96.38 83.505 97.14 ;
    RECT 26.71 95.62 26.88 96.38 ;
    RECT 26.88 95.53 27.16 96.47 ;
    RECT 27.16 95.62 27.32 96.38 ;
    RECT 27.8 95.62 28.02 96.38 ;
    RECT 28.5 95.62 28.72 96.38 ;
    RECT 29.2 95.62 30.815 96.38 ;
    RECT 31.295 95.62 31.515 96.38 ;
    RECT 31.995 95.62 32.21 96.38 ;
    RECT 32.69 95.62 32.91 96.38 ;
    RECT 33.39 95.62 33.61 96.38 ;
    RECT 34.09 95.62 34.31 96.38 ;
    RECT 34.79 95.62 35.005 96.38 ;
    RECT 35.485 95.62 36.405 96.38 ;
    RECT 36.885 95.62 37.105 96.38 ;
    RECT 37.585 95.62 37.8 96.38 ;
    RECT 38.28 95.62 38.5 96.38 ;
    RECT 38.98 95.62 39.2 96.38 ;
    RECT 39.68 95.62 39.895 96.38 ;
    RECT 40.375 95.62 40.595 96.38 ;
    RECT 41.075 95.62 41.995 96.38 ;
    RECT 42.475 95.62 42.69 96.38 ;
    RECT 43.17 95.62 43.39 96.38 ;
    RECT 43.87 95.62 44.09 96.38 ;
    RECT 44.57 95.62 44.79 96.38 ;
    RECT 45.27 95.62 45.485 96.38 ;
    RECT 45.965 95.62 46.185 96.38 ;
    RECT 46.665 95.62 47.58 96.38 ;
    RECT 48.06 95.62 48.28 96.38 ;
    RECT 48.76 95.62 48.98 96.38 ;
    RECT 49.46 95.62 49.68 96.38 ;
    RECT 50.16 95.62 50.375 96.38 ;
    RECT 50.855 95.62 51.775 96.38 ;
    RECT 52.255 95.62 53.17 96.38 ;
    RECT 53.65 95.62 53.87 96.38 ;
    RECT 54.35 95.62 54.57 96.38 ;
    RECT 55.05 95.62 55.265 96.38 ;
    RECT 55.745 95.62 55.965 96.38 ;
    RECT 56.445 95.62 56.665 96.38 ;
    RECT 57.145 95.62 58.06 96.38 ;
    RECT 58.54 95.62 59.46 96.38 ;
    RECT 59.94 95.62 60.16 96.38 ;
    RECT 60.64 95.62 60.855 96.38 ;
    RECT 61.335 95.62 61.555 96.38 ;
    RECT 62.035 95.62 62.25 96.38 ;
    RECT 62.73 95.62 63.65 96.38 ;
    RECT 64.13 95.62 64.345 96.38 ;
    RECT 64.825 95.62 65.045 96.38 ;
    RECT 65.525 95.62 65.745 96.38 ;
    RECT 66.225 95.62 66.445 96.38 ;
    RECT 66.925 95.62 67.14 96.38 ;
    RECT 67.62 95.62 67.84 96.38 ;
    RECT 68.32 95.62 69.235 96.38 ;
    RECT 69.715 95.62 69.935 96.38 ;
    RECT 70.415 95.62 70.635 96.38 ;
    RECT 71.115 95.62 71.335 96.38 ;
    RECT 71.815 95.62 72.035 96.38 ;
    RECT 72.515 95.62 72.735 96.38 ;
    RECT 73.215 95.62 73.435 96.38 ;
    RECT 73.915 95.62 74.835 96.38 ;
    RECT 75.315 95.62 75.535 96.38 ;
    RECT 76.015 95.62 76.225 96.38 ;
    RECT 76.705 95.62 76.92 96.38 ;
    RECT 77.4 95.62 77.62 96.38 ;
    RECT 78.1 95.62 78.32 96.38 ;
    RECT 78.8 95.62 79.02 96.38 ;
    RECT 79.5 95.62 81.115 96.38 ;
    RECT 81.595 95.62 81.815 96.38 ;
    RECT 82.295 95.62 82.515 96.38 ;
    RECT 82.995 95.62 83.055 96.38 ;
    RECT 83.055 95.53 83.335 96.47 ;
    RECT 83.335 95.62 83.505 96.38 ;
    RECT 26.71 94.86 26.88 95.62 ;
    RECT 26.88 94.77 27.16 95.71 ;
    RECT 27.16 94.86 27.32 95.62 ;
    RECT 27.8 94.86 28.02 95.62 ;
    RECT 28.5 94.86 28.72 95.62 ;
    RECT 29.2 94.86 30.815 95.62 ;
    RECT 31.295 94.86 31.515 95.62 ;
    RECT 31.995 94.86 32.21 95.62 ;
    RECT 32.69 94.86 32.91 95.62 ;
    RECT 33.39 94.86 33.61 95.62 ;
    RECT 34.09 94.86 34.31 95.62 ;
    RECT 34.79 94.86 35.005 95.62 ;
    RECT 35.485 94.86 36.405 95.62 ;
    RECT 36.885 94.86 37.105 95.62 ;
    RECT 37.585 94.86 37.8 95.62 ;
    RECT 38.28 94.86 38.5 95.62 ;
    RECT 38.98 94.86 39.2 95.62 ;
    RECT 39.68 94.86 39.895 95.62 ;
    RECT 40.375 94.86 40.595 95.62 ;
    RECT 41.075 94.86 41.995 95.62 ;
    RECT 42.475 94.86 42.69 95.62 ;
    RECT 43.17 94.86 43.39 95.62 ;
    RECT 43.87 94.86 44.09 95.62 ;
    RECT 44.57 94.86 44.79 95.62 ;
    RECT 45.27 94.86 45.485 95.62 ;
    RECT 45.965 94.86 46.185 95.62 ;
    RECT 46.665 94.86 47.58 95.62 ;
    RECT 48.06 94.86 48.28 95.62 ;
    RECT 48.76 94.86 48.98 95.62 ;
    RECT 49.46 94.86 49.68 95.62 ;
    RECT 50.16 94.86 50.375 95.62 ;
    RECT 50.855 94.86 51.775 95.62 ;
    RECT 52.255 94.86 53.17 95.62 ;
    RECT 53.65 94.86 53.87 95.62 ;
    RECT 54.35 94.86 54.57 95.62 ;
    RECT 55.05 94.86 55.265 95.62 ;
    RECT 55.745 94.86 55.965 95.62 ;
    RECT 56.445 94.86 56.665 95.62 ;
    RECT 57.145 94.86 58.06 95.62 ;
    RECT 58.54 94.86 59.46 95.62 ;
    RECT 59.94 94.86 60.16 95.62 ;
    RECT 60.64 94.86 60.855 95.62 ;
    RECT 61.335 94.86 61.555 95.62 ;
    RECT 62.035 94.86 62.25 95.62 ;
    RECT 62.73 94.86 63.65 95.62 ;
    RECT 64.13 94.86 64.345 95.62 ;
    RECT 64.825 94.86 65.045 95.62 ;
    RECT 65.525 94.86 65.745 95.62 ;
    RECT 66.225 94.86 66.445 95.62 ;
    RECT 66.925 94.86 67.14 95.62 ;
    RECT 67.62 94.86 67.84 95.62 ;
    RECT 68.32 94.86 69.235 95.62 ;
    RECT 69.715 94.86 69.935 95.62 ;
    RECT 70.415 94.86 70.635 95.62 ;
    RECT 71.115 94.86 71.335 95.62 ;
    RECT 71.815 94.86 72.035 95.62 ;
    RECT 72.515 94.86 72.735 95.62 ;
    RECT 73.215 94.86 73.435 95.62 ;
    RECT 73.915 94.86 74.835 95.62 ;
    RECT 75.315 94.86 75.535 95.62 ;
    RECT 76.015 94.86 76.225 95.62 ;
    RECT 76.705 94.86 76.92 95.62 ;
    RECT 77.4 94.86 77.62 95.62 ;
    RECT 78.1 94.86 78.32 95.62 ;
    RECT 78.8 94.86 79.02 95.62 ;
    RECT 79.5 94.86 81.115 95.62 ;
    RECT 81.595 94.86 81.815 95.62 ;
    RECT 82.295 94.86 82.515 95.62 ;
    RECT 82.995 94.86 83.055 95.62 ;
    RECT 83.055 94.77 83.335 95.71 ;
    RECT 83.335 94.86 83.505 95.62 ;
    RECT 26.71 94.1 26.88 94.86 ;
    RECT 26.88 94.01 27.16 94.95 ;
    RECT 27.16 94.1 27.32 94.86 ;
    RECT 27.8 94.1 28.02 94.86 ;
    RECT 28.5 94.1 28.72 94.86 ;
    RECT 29.2 94.1 30.815 94.86 ;
    RECT 31.295 94.1 31.515 94.86 ;
    RECT 31.995 94.1 32.21 94.86 ;
    RECT 32.69 94.1 32.91 94.86 ;
    RECT 33.39 94.1 33.61 94.86 ;
    RECT 34.09 94.1 34.31 94.86 ;
    RECT 34.79 94.1 35.005 94.86 ;
    RECT 35.485 94.1 36.405 94.86 ;
    RECT 36.885 94.1 37.105 94.86 ;
    RECT 37.585 94.1 37.8 94.86 ;
    RECT 38.28 94.1 38.5 94.86 ;
    RECT 38.98 94.1 39.2 94.86 ;
    RECT 39.68 94.1 39.895 94.86 ;
    RECT 40.375 94.1 40.595 94.86 ;
    RECT 41.075 94.1 41.995 94.86 ;
    RECT 42.475 94.1 42.69 94.86 ;
    RECT 43.17 94.1 43.39 94.86 ;
    RECT 43.87 94.1 44.09 94.86 ;
    RECT 44.57 94.1 44.79 94.86 ;
    RECT 45.27 94.1 45.485 94.86 ;
    RECT 45.965 94.1 46.185 94.86 ;
    RECT 46.665 94.1 47.58 94.86 ;
    RECT 48.06 94.1 48.28 94.86 ;
    RECT 48.76 94.1 48.98 94.86 ;
    RECT 49.46 94.1 49.68 94.86 ;
    RECT 50.16 94.1 50.375 94.86 ;
    RECT 50.855 94.1 51.775 94.86 ;
    RECT 52.255 94.1 53.17 94.86 ;
    RECT 53.65 94.1 53.87 94.86 ;
    RECT 54.35 94.1 54.57 94.86 ;
    RECT 55.05 94.1 55.265 94.86 ;
    RECT 55.745 94.1 55.965 94.86 ;
    RECT 56.445 94.1 56.665 94.86 ;
    RECT 57.145 94.1 58.06 94.86 ;
    RECT 58.54 94.1 59.46 94.86 ;
    RECT 59.94 94.1 60.16 94.86 ;
    RECT 60.64 94.1 60.855 94.86 ;
    RECT 61.335 94.1 61.555 94.86 ;
    RECT 62.035 94.1 62.25 94.86 ;
    RECT 62.73 94.1 63.65 94.86 ;
    RECT 64.13 94.1 64.345 94.86 ;
    RECT 64.825 94.1 65.045 94.86 ;
    RECT 65.525 94.1 65.745 94.86 ;
    RECT 66.225 94.1 66.445 94.86 ;
    RECT 66.925 94.1 67.14 94.86 ;
    RECT 67.62 94.1 67.84 94.86 ;
    RECT 68.32 94.1 69.235 94.86 ;
    RECT 69.715 94.1 69.935 94.86 ;
    RECT 70.415 94.1 70.635 94.86 ;
    RECT 71.115 94.1 71.335 94.86 ;
    RECT 71.815 94.1 72.035 94.86 ;
    RECT 72.515 94.1 72.735 94.86 ;
    RECT 73.215 94.1 73.435 94.86 ;
    RECT 73.915 94.1 74.835 94.86 ;
    RECT 75.315 94.1 75.535 94.86 ;
    RECT 76.015 94.1 76.225 94.86 ;
    RECT 76.705 94.1 76.92 94.86 ;
    RECT 77.4 94.1 77.62 94.86 ;
    RECT 78.1 94.1 78.32 94.86 ;
    RECT 78.8 94.1 79.02 94.86 ;
    RECT 79.5 94.1 81.115 94.86 ;
    RECT 81.595 94.1 81.815 94.86 ;
    RECT 82.295 94.1 82.515 94.86 ;
    RECT 82.995 94.1 83.055 94.86 ;
    RECT 83.055 94.01 83.335 94.95 ;
    RECT 83.335 94.1 83.505 94.86 ;
    RECT 26.71 93.34 26.88 94.1 ;
    RECT 26.88 93.25 27.16 94.19 ;
    RECT 27.16 93.34 27.32 94.1 ;
    RECT 27.8 93.34 28.02 94.1 ;
    RECT 28.5 93.34 28.72 94.1 ;
    RECT 29.2 93.34 30.815 94.1 ;
    RECT 31.295 93.34 31.515 94.1 ;
    RECT 31.995 93.34 32.21 94.1 ;
    RECT 32.69 93.34 32.91 94.1 ;
    RECT 33.39 93.34 33.61 94.1 ;
    RECT 34.09 93.34 34.31 94.1 ;
    RECT 34.79 93.34 35.005 94.1 ;
    RECT 35.485 93.34 36.405 94.1 ;
    RECT 36.885 93.34 37.105 94.1 ;
    RECT 37.585 93.34 37.8 94.1 ;
    RECT 38.28 93.34 38.5 94.1 ;
    RECT 38.98 93.34 39.2 94.1 ;
    RECT 39.68 93.34 39.895 94.1 ;
    RECT 40.375 93.34 40.595 94.1 ;
    RECT 41.075 93.34 41.995 94.1 ;
    RECT 42.475 93.34 42.69 94.1 ;
    RECT 43.17 93.34 43.39 94.1 ;
    RECT 43.87 93.34 44.09 94.1 ;
    RECT 44.57 93.34 44.79 94.1 ;
    RECT 45.27 93.34 45.485 94.1 ;
    RECT 45.965 93.34 46.185 94.1 ;
    RECT 46.665 93.34 47.58 94.1 ;
    RECT 48.06 93.34 48.28 94.1 ;
    RECT 48.76 93.34 48.98 94.1 ;
    RECT 49.46 93.34 49.68 94.1 ;
    RECT 50.16 93.34 50.375 94.1 ;
    RECT 50.855 93.34 51.775 94.1 ;
    RECT 52.255 93.34 53.17 94.1 ;
    RECT 53.65 93.34 53.87 94.1 ;
    RECT 54.35 93.34 54.57 94.1 ;
    RECT 55.05 93.34 55.265 94.1 ;
    RECT 55.745 93.34 55.965 94.1 ;
    RECT 56.445 93.34 56.665 94.1 ;
    RECT 57.145 93.34 58.06 94.1 ;
    RECT 58.54 93.34 59.46 94.1 ;
    RECT 59.94 93.34 60.16 94.1 ;
    RECT 60.64 93.34 60.855 94.1 ;
    RECT 61.335 93.34 61.555 94.1 ;
    RECT 62.035 93.34 62.25 94.1 ;
    RECT 62.73 93.34 63.65 94.1 ;
    RECT 64.13 93.34 64.345 94.1 ;
    RECT 64.825 93.34 65.045 94.1 ;
    RECT 65.525 93.34 65.745 94.1 ;
    RECT 66.225 93.34 66.445 94.1 ;
    RECT 66.925 93.34 67.14 94.1 ;
    RECT 67.62 93.34 67.84 94.1 ;
    RECT 68.32 93.34 69.235 94.1 ;
    RECT 69.715 93.34 69.935 94.1 ;
    RECT 70.415 93.34 70.635 94.1 ;
    RECT 71.115 93.34 71.335 94.1 ;
    RECT 71.815 93.34 72.035 94.1 ;
    RECT 72.515 93.34 72.735 94.1 ;
    RECT 73.215 93.34 73.435 94.1 ;
    RECT 73.915 93.34 74.835 94.1 ;
    RECT 75.315 93.34 75.535 94.1 ;
    RECT 76.015 93.34 76.225 94.1 ;
    RECT 76.705 93.34 76.92 94.1 ;
    RECT 77.4 93.34 77.62 94.1 ;
    RECT 78.1 93.34 78.32 94.1 ;
    RECT 78.8 93.34 79.02 94.1 ;
    RECT 79.5 93.34 81.115 94.1 ;
    RECT 81.595 93.34 81.815 94.1 ;
    RECT 82.295 93.34 82.515 94.1 ;
    RECT 82.995 93.34 83.055 94.1 ;
    RECT 83.055 93.25 83.335 94.19 ;
    RECT 83.335 93.34 83.505 94.1 ;
    RECT 26.71 92.58 26.88 93.34 ;
    RECT 26.88 92.49 27.16 93.43 ;
    RECT 27.16 92.58 27.32 93.34 ;
    RECT 27.8 92.58 28.02 93.34 ;
    RECT 28.5 92.58 28.72 93.34 ;
    RECT 29.2 92.58 30.815 93.34 ;
    RECT 31.295 92.58 31.515 93.34 ;
    RECT 31.995 92.58 32.21 93.34 ;
    RECT 32.69 92.58 32.91 93.34 ;
    RECT 33.39 92.58 33.61 93.34 ;
    RECT 34.09 92.58 34.31 93.34 ;
    RECT 34.79 92.58 35.005 93.34 ;
    RECT 35.485 92.58 36.405 93.34 ;
    RECT 36.885 92.58 37.105 93.34 ;
    RECT 37.585 92.58 37.8 93.34 ;
    RECT 38.28 92.58 38.5 93.34 ;
    RECT 38.98 92.58 39.2 93.34 ;
    RECT 39.68 92.58 39.895 93.34 ;
    RECT 40.375 92.58 40.595 93.34 ;
    RECT 41.075 92.58 41.995 93.34 ;
    RECT 42.475 92.58 42.69 93.34 ;
    RECT 43.17 92.58 43.39 93.34 ;
    RECT 43.87 92.58 44.09 93.34 ;
    RECT 44.57 92.58 44.79 93.34 ;
    RECT 45.27 92.58 45.485 93.34 ;
    RECT 45.965 92.58 46.185 93.34 ;
    RECT 46.665 92.58 47.58 93.34 ;
    RECT 48.06 92.58 48.28 93.34 ;
    RECT 48.76 92.58 48.98 93.34 ;
    RECT 49.46 92.58 49.68 93.34 ;
    RECT 50.16 92.58 50.375 93.34 ;
    RECT 50.855 92.58 51.775 93.34 ;
    RECT 52.255 92.58 53.17 93.34 ;
    RECT 53.65 92.58 53.87 93.34 ;
    RECT 54.35 92.58 54.57 93.34 ;
    RECT 55.05 92.58 55.265 93.34 ;
    RECT 55.745 92.58 55.965 93.34 ;
    RECT 56.445 92.58 56.665 93.34 ;
    RECT 57.145 92.58 58.06 93.34 ;
    RECT 58.54 92.58 59.46 93.34 ;
    RECT 59.94 92.58 60.16 93.34 ;
    RECT 60.64 92.58 60.855 93.34 ;
    RECT 61.335 92.58 61.555 93.34 ;
    RECT 62.035 92.58 62.25 93.34 ;
    RECT 62.73 92.58 63.65 93.34 ;
    RECT 64.13 92.58 64.345 93.34 ;
    RECT 64.825 92.58 65.045 93.34 ;
    RECT 65.525 92.58 65.745 93.34 ;
    RECT 66.225 92.58 66.445 93.34 ;
    RECT 66.925 92.58 67.14 93.34 ;
    RECT 67.62 92.58 67.84 93.34 ;
    RECT 68.32 92.58 69.235 93.34 ;
    RECT 69.715 92.58 69.935 93.34 ;
    RECT 70.415 92.58 70.635 93.34 ;
    RECT 71.115 92.58 71.335 93.34 ;
    RECT 71.815 92.58 72.035 93.34 ;
    RECT 72.515 92.58 72.735 93.34 ;
    RECT 73.215 92.58 73.435 93.34 ;
    RECT 73.915 92.58 74.835 93.34 ;
    RECT 75.315 92.58 75.535 93.34 ;
    RECT 76.015 92.58 76.225 93.34 ;
    RECT 76.705 92.58 76.92 93.34 ;
    RECT 77.4 92.58 77.62 93.34 ;
    RECT 78.1 92.58 78.32 93.34 ;
    RECT 78.8 92.58 79.02 93.34 ;
    RECT 79.5 92.58 81.115 93.34 ;
    RECT 81.595 92.58 81.815 93.34 ;
    RECT 82.295 92.58 82.515 93.34 ;
    RECT 82.995 92.58 83.055 93.34 ;
    RECT 83.055 92.49 83.335 93.43 ;
    RECT 83.335 92.58 83.505 93.34 ;
    RECT 26.71 91.82 26.88 92.58 ;
    RECT 26.88 91.73 27.16 92.67 ;
    RECT 27.16 91.82 27.32 92.58 ;
    RECT 27.8 91.82 28.02 92.58 ;
    RECT 28.5 91.82 28.72 92.58 ;
    RECT 29.2 91.82 30.815 92.58 ;
    RECT 31.295 91.82 31.515 92.58 ;
    RECT 31.995 91.82 32.21 92.58 ;
    RECT 32.69 91.82 32.91 92.58 ;
    RECT 33.39 91.82 33.61 92.58 ;
    RECT 34.09 91.82 34.31 92.58 ;
    RECT 34.79 91.82 35.005 92.58 ;
    RECT 35.485 91.82 36.405 92.58 ;
    RECT 36.885 91.82 37.105 92.58 ;
    RECT 37.585 91.82 37.8 92.58 ;
    RECT 38.28 91.82 38.5 92.58 ;
    RECT 38.98 91.82 39.2 92.58 ;
    RECT 39.68 91.82 39.895 92.58 ;
    RECT 40.375 91.82 40.595 92.58 ;
    RECT 41.075 91.82 41.995 92.58 ;
    RECT 42.475 91.82 42.69 92.58 ;
    RECT 43.17 91.82 43.39 92.58 ;
    RECT 43.87 91.82 44.09 92.58 ;
    RECT 44.57 91.82 44.79 92.58 ;
    RECT 45.27 91.82 45.485 92.58 ;
    RECT 45.965 91.82 46.185 92.58 ;
    RECT 46.665 91.82 47.58 92.58 ;
    RECT 48.06 91.82 48.28 92.58 ;
    RECT 48.76 91.82 48.98 92.58 ;
    RECT 49.46 91.82 49.68 92.58 ;
    RECT 50.16 91.82 50.375 92.58 ;
    RECT 50.855 91.82 51.775 92.58 ;
    RECT 52.255 91.82 53.17 92.58 ;
    RECT 53.65 91.82 53.87 92.58 ;
    RECT 54.35 91.82 54.57 92.58 ;
    RECT 55.05 91.82 55.265 92.58 ;
    RECT 55.745 91.82 55.965 92.58 ;
    RECT 56.445 91.82 56.665 92.58 ;
    RECT 57.145 91.82 58.06 92.58 ;
    RECT 58.54 91.82 59.46 92.58 ;
    RECT 59.94 91.82 60.16 92.58 ;
    RECT 60.64 91.82 60.855 92.58 ;
    RECT 61.335 91.82 61.555 92.58 ;
    RECT 62.035 91.82 62.25 92.58 ;
    RECT 62.73 91.82 63.65 92.58 ;
    RECT 64.13 91.82 64.345 92.58 ;
    RECT 64.825 91.82 65.045 92.58 ;
    RECT 65.525 91.82 65.745 92.58 ;
    RECT 66.225 91.82 66.445 92.58 ;
    RECT 66.925 91.82 67.14 92.58 ;
    RECT 67.62 91.82 67.84 92.58 ;
    RECT 68.32 91.82 69.235 92.58 ;
    RECT 69.715 91.82 69.935 92.58 ;
    RECT 70.415 91.82 70.635 92.58 ;
    RECT 71.115 91.82 71.335 92.58 ;
    RECT 71.815 91.82 72.035 92.58 ;
    RECT 72.515 91.82 72.735 92.58 ;
    RECT 73.215 91.82 73.435 92.58 ;
    RECT 73.915 91.82 74.835 92.58 ;
    RECT 75.315 91.82 75.535 92.58 ;
    RECT 76.015 91.82 76.225 92.58 ;
    RECT 76.705 91.82 76.92 92.58 ;
    RECT 77.4 91.82 77.62 92.58 ;
    RECT 78.1 91.82 78.32 92.58 ;
    RECT 78.8 91.82 79.02 92.58 ;
    RECT 79.5 91.82 81.115 92.58 ;
    RECT 81.595 91.82 81.815 92.58 ;
    RECT 82.295 91.82 82.515 92.58 ;
    RECT 82.995 91.82 83.055 92.58 ;
    RECT 83.055 91.73 83.335 92.67 ;
    RECT 83.335 91.82 83.505 92.58 ;
    RECT 26.71 91.06 26.88 91.82 ;
    RECT 26.88 90.97 27.16 91.91 ;
    RECT 27.16 91.06 27.32 91.82 ;
    RECT 27.8 91.06 28.02 91.82 ;
    RECT 28.5 91.06 28.72 91.82 ;
    RECT 29.2 91.06 30.815 91.82 ;
    RECT 31.295 91.06 31.515 91.82 ;
    RECT 31.995 91.06 32.21 91.82 ;
    RECT 32.69 91.06 32.91 91.82 ;
    RECT 33.39 91.06 33.61 91.82 ;
    RECT 34.09 91.06 34.31 91.82 ;
    RECT 34.79 91.06 35.005 91.82 ;
    RECT 35.485 91.06 36.405 91.82 ;
    RECT 36.885 91.06 37.105 91.82 ;
    RECT 37.585 91.06 37.8 91.82 ;
    RECT 38.28 91.06 38.5 91.82 ;
    RECT 38.98 91.06 39.2 91.82 ;
    RECT 39.68 91.06 39.895 91.82 ;
    RECT 40.375 91.06 40.595 91.82 ;
    RECT 41.075 91.06 41.995 91.82 ;
    RECT 42.475 91.06 42.69 91.82 ;
    RECT 43.17 91.06 43.39 91.82 ;
    RECT 43.87 91.06 44.09 91.82 ;
    RECT 44.57 91.06 44.79 91.82 ;
    RECT 45.27 91.06 45.485 91.82 ;
    RECT 45.965 91.06 46.185 91.82 ;
    RECT 46.665 91.06 47.58 91.82 ;
    RECT 48.06 91.06 48.28 91.82 ;
    RECT 48.76 91.06 48.98 91.82 ;
    RECT 49.46 91.06 49.68 91.82 ;
    RECT 50.16 91.06 50.375 91.82 ;
    RECT 50.855 91.06 51.775 91.82 ;
    RECT 52.255 91.06 53.17 91.82 ;
    RECT 53.65 91.06 53.87 91.82 ;
    RECT 54.35 91.06 54.57 91.82 ;
    RECT 55.05 91.06 55.265 91.82 ;
    RECT 55.745 91.06 55.965 91.82 ;
    RECT 56.445 91.06 56.665 91.82 ;
    RECT 57.145 91.06 58.06 91.82 ;
    RECT 58.54 91.06 59.46 91.82 ;
    RECT 59.94 91.06 60.16 91.82 ;
    RECT 60.64 91.06 60.855 91.82 ;
    RECT 61.335 91.06 61.555 91.82 ;
    RECT 62.035 91.06 62.25 91.82 ;
    RECT 62.73 91.06 63.65 91.82 ;
    RECT 64.13 91.06 64.345 91.82 ;
    RECT 64.825 91.06 65.045 91.82 ;
    RECT 65.525 91.06 65.745 91.82 ;
    RECT 66.225 91.06 66.445 91.82 ;
    RECT 66.925 91.06 67.14 91.82 ;
    RECT 67.62 91.06 67.84 91.82 ;
    RECT 68.32 91.06 69.235 91.82 ;
    RECT 69.715 91.06 69.935 91.82 ;
    RECT 70.415 91.06 70.635 91.82 ;
    RECT 71.115 91.06 71.335 91.82 ;
    RECT 71.815 91.06 72.035 91.82 ;
    RECT 72.515 91.06 72.735 91.82 ;
    RECT 73.215 91.06 73.435 91.82 ;
    RECT 73.915 91.06 74.835 91.82 ;
    RECT 75.315 91.06 75.535 91.82 ;
    RECT 76.015 91.06 76.225 91.82 ;
    RECT 76.705 91.06 76.92 91.82 ;
    RECT 77.4 91.06 77.62 91.82 ;
    RECT 78.1 91.06 78.32 91.82 ;
    RECT 78.8 91.06 79.02 91.82 ;
    RECT 79.5 91.06 81.115 91.82 ;
    RECT 81.595 91.06 81.815 91.82 ;
    RECT 82.295 91.06 82.515 91.82 ;
    RECT 82.995 91.06 83.055 91.82 ;
    RECT 83.055 90.97 83.335 91.91 ;
    RECT 83.335 91.06 83.505 91.82 ;
    RECT 26.71 90.3 26.88 91.06 ;
    RECT 26.88 90.21 27.16 91.15 ;
    RECT 27.16 90.3 27.32 91.06 ;
    RECT 27.8 90.3 28.02 91.06 ;
    RECT 28.5 90.3 28.72 91.06 ;
    RECT 29.2 90.3 30.815 91.06 ;
    RECT 31.295 90.3 31.515 91.06 ;
    RECT 31.995 90.3 32.21 91.06 ;
    RECT 32.69 90.3 32.91 91.06 ;
    RECT 33.39 90.3 33.61 91.06 ;
    RECT 34.09 90.3 34.31 91.06 ;
    RECT 34.79 90.3 35.005 91.06 ;
    RECT 35.485 90.3 36.405 91.06 ;
    RECT 36.885 90.3 37.105 91.06 ;
    RECT 37.585 90.3 37.8 91.06 ;
    RECT 38.28 90.3 38.5 91.06 ;
    RECT 38.98 90.3 39.2 91.06 ;
    RECT 39.68 90.3 39.895 91.06 ;
    RECT 40.375 90.3 40.595 91.06 ;
    RECT 41.075 90.3 41.995 91.06 ;
    RECT 42.475 90.3 42.69 91.06 ;
    RECT 43.17 90.3 43.39 91.06 ;
    RECT 43.87 90.3 44.09 91.06 ;
    RECT 44.57 90.3 44.79 91.06 ;
    RECT 45.27 90.3 45.485 91.06 ;
    RECT 45.965 90.3 46.185 91.06 ;
    RECT 46.665 90.3 47.58 91.06 ;
    RECT 48.06 90.3 48.28 91.06 ;
    RECT 48.76 90.3 48.98 91.06 ;
    RECT 49.46 90.3 49.68 91.06 ;
    RECT 50.16 90.3 50.375 91.06 ;
    RECT 50.855 90.3 51.775 91.06 ;
    RECT 52.255 90.3 53.17 91.06 ;
    RECT 53.65 90.3 53.87 91.06 ;
    RECT 54.35 90.3 54.57 91.06 ;
    RECT 55.05 90.3 55.265 91.06 ;
    RECT 55.745 90.3 55.965 91.06 ;
    RECT 56.445 90.3 56.665 91.06 ;
    RECT 57.145 90.3 58.06 91.06 ;
    RECT 58.54 90.3 59.46 91.06 ;
    RECT 59.94 90.3 60.16 91.06 ;
    RECT 60.64 90.3 60.855 91.06 ;
    RECT 61.335 90.3 61.555 91.06 ;
    RECT 62.035 90.3 62.25 91.06 ;
    RECT 62.73 90.3 63.65 91.06 ;
    RECT 64.13 90.3 64.345 91.06 ;
    RECT 64.825 90.3 65.045 91.06 ;
    RECT 65.525 90.3 65.745 91.06 ;
    RECT 66.225 90.3 66.445 91.06 ;
    RECT 66.925 90.3 67.14 91.06 ;
    RECT 67.62 90.3 67.84 91.06 ;
    RECT 68.32 90.3 69.235 91.06 ;
    RECT 69.715 90.3 69.935 91.06 ;
    RECT 70.415 90.3 70.635 91.06 ;
    RECT 71.115 90.3 71.335 91.06 ;
    RECT 71.815 90.3 72.035 91.06 ;
    RECT 72.515 90.3 72.735 91.06 ;
    RECT 73.215 90.3 73.435 91.06 ;
    RECT 73.915 90.3 74.835 91.06 ;
    RECT 75.315 90.3 75.535 91.06 ;
    RECT 76.015 90.3 76.225 91.06 ;
    RECT 76.705 90.3 76.92 91.06 ;
    RECT 77.4 90.3 77.62 91.06 ;
    RECT 78.1 90.3 78.32 91.06 ;
    RECT 78.8 90.3 79.02 91.06 ;
    RECT 79.5 90.3 81.115 91.06 ;
    RECT 81.595 90.3 81.815 91.06 ;
    RECT 82.295 90.3 82.515 91.06 ;
    RECT 82.995 90.3 83.055 91.06 ;
    RECT 83.055 90.21 83.335 91.15 ;
    RECT 83.335 90.3 83.505 91.06 ;
    RECT 26.71 89.54 26.88 90.3 ;
    RECT 26.88 89.45 27.16 90.39 ;
    RECT 27.16 89.54 27.32 90.3 ;
    RECT 27.8 89.54 28.02 90.3 ;
    RECT 28.5 89.54 28.72 90.3 ;
    RECT 29.2 89.54 30.815 90.3 ;
    RECT 31.295 89.54 31.515 90.3 ;
    RECT 31.995 89.54 32.21 90.3 ;
    RECT 32.69 89.54 32.91 90.3 ;
    RECT 33.39 89.54 33.61 90.3 ;
    RECT 34.09 89.54 34.31 90.3 ;
    RECT 34.79 89.54 35.005 90.3 ;
    RECT 35.485 89.54 36.405 90.3 ;
    RECT 36.885 89.54 37.105 90.3 ;
    RECT 37.585 89.54 37.8 90.3 ;
    RECT 38.28 89.54 38.5 90.3 ;
    RECT 38.98 89.54 39.2 90.3 ;
    RECT 39.68 89.54 39.895 90.3 ;
    RECT 40.375 89.54 40.595 90.3 ;
    RECT 41.075 89.54 41.995 90.3 ;
    RECT 42.475 89.54 42.69 90.3 ;
    RECT 43.17 89.54 43.39 90.3 ;
    RECT 43.87 89.54 44.09 90.3 ;
    RECT 44.57 89.54 44.79 90.3 ;
    RECT 45.27 89.54 45.485 90.3 ;
    RECT 45.965 89.54 46.185 90.3 ;
    RECT 46.665 89.54 47.58 90.3 ;
    RECT 48.06 89.54 48.28 90.3 ;
    RECT 48.76 89.54 48.98 90.3 ;
    RECT 49.46 89.54 49.68 90.3 ;
    RECT 50.16 89.54 50.375 90.3 ;
    RECT 50.855 89.54 51.775 90.3 ;
    RECT 52.255 89.54 53.17 90.3 ;
    RECT 53.65 89.54 53.87 90.3 ;
    RECT 54.35 89.54 54.57 90.3 ;
    RECT 55.05 89.54 55.265 90.3 ;
    RECT 55.745 89.54 55.965 90.3 ;
    RECT 56.445 89.54 56.665 90.3 ;
    RECT 57.145 89.54 58.06 90.3 ;
    RECT 58.54 89.54 59.46 90.3 ;
    RECT 59.94 89.54 60.16 90.3 ;
    RECT 60.64 89.54 60.855 90.3 ;
    RECT 61.335 89.54 61.555 90.3 ;
    RECT 62.035 89.54 62.25 90.3 ;
    RECT 62.73 89.54 63.65 90.3 ;
    RECT 64.13 89.54 64.345 90.3 ;
    RECT 64.825 89.54 65.045 90.3 ;
    RECT 65.525 89.54 65.745 90.3 ;
    RECT 66.225 89.54 66.445 90.3 ;
    RECT 66.925 89.54 67.14 90.3 ;
    RECT 67.62 89.54 67.84 90.3 ;
    RECT 68.32 89.54 69.235 90.3 ;
    RECT 69.715 89.54 69.935 90.3 ;
    RECT 70.415 89.54 70.635 90.3 ;
    RECT 71.115 89.54 71.335 90.3 ;
    RECT 71.815 89.54 72.035 90.3 ;
    RECT 72.515 89.54 72.735 90.3 ;
    RECT 73.215 89.54 73.435 90.3 ;
    RECT 73.915 89.54 74.835 90.3 ;
    RECT 75.315 89.54 75.535 90.3 ;
    RECT 76.015 89.54 76.225 90.3 ;
    RECT 76.705 89.54 76.92 90.3 ;
    RECT 77.4 89.54 77.62 90.3 ;
    RECT 78.1 89.54 78.32 90.3 ;
    RECT 78.8 89.54 79.02 90.3 ;
    RECT 79.5 89.54 81.115 90.3 ;
    RECT 81.595 89.54 81.815 90.3 ;
    RECT 82.295 89.54 82.515 90.3 ;
    RECT 82.995 89.54 83.055 90.3 ;
    RECT 83.055 89.45 83.335 90.39 ;
    RECT 83.335 89.54 83.505 90.3 ;
    RECT 26.71 88.78 26.88 89.54 ;
    RECT 26.88 88.69 27.16 89.63 ;
    RECT 27.16 88.78 27.32 89.54 ;
    RECT 27.8 88.78 28.02 89.54 ;
    RECT 28.5 88.78 28.72 89.54 ;
    RECT 29.2 88.78 30.815 89.54 ;
    RECT 31.295 88.78 31.515 89.54 ;
    RECT 31.995 88.78 32.21 89.54 ;
    RECT 32.69 88.78 32.91 89.54 ;
    RECT 33.39 88.78 33.61 89.54 ;
    RECT 34.09 88.78 34.31 89.54 ;
    RECT 34.79 88.78 35.005 89.54 ;
    RECT 35.485 88.78 36.405 89.54 ;
    RECT 36.885 88.78 37.105 89.54 ;
    RECT 37.585 88.78 37.8 89.54 ;
    RECT 38.28 88.78 38.5 89.54 ;
    RECT 38.98 88.78 39.2 89.54 ;
    RECT 39.68 88.78 39.895 89.54 ;
    RECT 40.375 88.78 40.595 89.54 ;
    RECT 41.075 88.78 41.995 89.54 ;
    RECT 42.475 88.78 42.69 89.54 ;
    RECT 43.17 88.78 43.39 89.54 ;
    RECT 43.87 88.78 44.09 89.54 ;
    RECT 44.57 88.78 44.79 89.54 ;
    RECT 45.27 88.78 45.485 89.54 ;
    RECT 45.965 88.78 46.185 89.54 ;
    RECT 46.665 88.78 47.58 89.54 ;
    RECT 48.06 88.78 48.28 89.54 ;
    RECT 48.76 88.78 48.98 89.54 ;
    RECT 49.46 88.78 49.68 89.54 ;
    RECT 50.16 88.78 50.375 89.54 ;
    RECT 50.855 88.78 51.775 89.54 ;
    RECT 52.255 88.78 53.17 89.54 ;
    RECT 53.65 88.78 53.87 89.54 ;
    RECT 54.35 88.78 54.57 89.54 ;
    RECT 55.05 88.78 55.265 89.54 ;
    RECT 55.745 88.78 55.965 89.54 ;
    RECT 56.445 88.78 56.665 89.54 ;
    RECT 57.145 88.78 58.06 89.54 ;
    RECT 58.54 88.78 59.46 89.54 ;
    RECT 59.94 88.78 60.16 89.54 ;
    RECT 60.64 88.78 60.855 89.54 ;
    RECT 61.335 88.78 61.555 89.54 ;
    RECT 62.035 88.78 62.25 89.54 ;
    RECT 62.73 88.78 63.65 89.54 ;
    RECT 64.13 88.78 64.345 89.54 ;
    RECT 64.825 88.78 65.045 89.54 ;
    RECT 65.525 88.78 65.745 89.54 ;
    RECT 66.225 88.78 66.445 89.54 ;
    RECT 66.925 88.78 67.14 89.54 ;
    RECT 67.62 88.78 67.84 89.54 ;
    RECT 68.32 88.78 69.235 89.54 ;
    RECT 69.715 88.78 69.935 89.54 ;
    RECT 70.415 88.78 70.635 89.54 ;
    RECT 71.115 88.78 71.335 89.54 ;
    RECT 71.815 88.78 72.035 89.54 ;
    RECT 72.515 88.78 72.735 89.54 ;
    RECT 73.215 88.78 73.435 89.54 ;
    RECT 73.915 88.78 74.835 89.54 ;
    RECT 75.315 88.78 75.535 89.54 ;
    RECT 76.015 88.78 76.225 89.54 ;
    RECT 76.705 88.78 76.92 89.54 ;
    RECT 77.4 88.78 77.62 89.54 ;
    RECT 78.1 88.78 78.32 89.54 ;
    RECT 78.8 88.78 79.02 89.54 ;
    RECT 79.5 88.78 81.115 89.54 ;
    RECT 81.595 88.78 81.815 89.54 ;
    RECT 82.295 88.78 82.515 89.54 ;
    RECT 82.995 88.78 83.055 89.54 ;
    RECT 83.055 88.69 83.335 89.63 ;
    RECT 83.335 88.78 83.505 89.54 ;
    RECT 26.71 88.02 26.88 88.78 ;
    RECT 26.88 87.93 27.16 88.87 ;
    RECT 27.16 88.02 27.32 88.78 ;
    RECT 27.8 88.02 28.02 88.78 ;
    RECT 28.5 88.02 28.72 88.78 ;
    RECT 29.2 88.02 30.815 88.78 ;
    RECT 31.295 88.02 31.515 88.78 ;
    RECT 31.995 88.02 32.21 88.78 ;
    RECT 32.69 88.02 32.91 88.78 ;
    RECT 33.39 88.02 33.61 88.78 ;
    RECT 34.09 88.02 34.31 88.78 ;
    RECT 34.79 88.02 35.005 88.78 ;
    RECT 35.485 88.02 36.405 88.78 ;
    RECT 36.885 88.02 37.105 88.78 ;
    RECT 37.585 88.02 37.8 88.78 ;
    RECT 38.28 88.02 38.5 88.78 ;
    RECT 38.98 88.02 39.2 88.78 ;
    RECT 39.68 88.02 39.895 88.78 ;
    RECT 40.375 88.02 40.595 88.78 ;
    RECT 41.075 88.02 41.995 88.78 ;
    RECT 42.475 88.02 42.69 88.78 ;
    RECT 43.17 88.02 43.39 88.78 ;
    RECT 43.87 88.02 44.09 88.78 ;
    RECT 44.57 88.02 44.79 88.78 ;
    RECT 45.27 88.02 45.485 88.78 ;
    RECT 45.965 88.02 46.185 88.78 ;
    RECT 46.665 88.02 47.58 88.78 ;
    RECT 48.06 88.02 48.28 88.78 ;
    RECT 48.76 88.02 48.98 88.78 ;
    RECT 49.46 88.02 49.68 88.78 ;
    RECT 50.16 88.02 50.375 88.78 ;
    RECT 50.855 88.02 51.775 88.78 ;
    RECT 52.255 88.02 53.17 88.78 ;
    RECT 53.65 88.02 53.87 88.78 ;
    RECT 54.35 88.02 54.57 88.78 ;
    RECT 55.05 88.02 55.265 88.78 ;
    RECT 55.745 88.02 55.965 88.78 ;
    RECT 56.445 88.02 56.665 88.78 ;
    RECT 57.145 88.02 58.06 88.78 ;
    RECT 58.54 88.02 59.46 88.78 ;
    RECT 59.94 88.02 60.16 88.78 ;
    RECT 60.64 88.02 60.855 88.78 ;
    RECT 61.335 88.02 61.555 88.78 ;
    RECT 62.035 88.02 62.25 88.78 ;
    RECT 62.73 88.02 63.65 88.78 ;
    RECT 64.13 88.02 64.345 88.78 ;
    RECT 64.825 88.02 65.045 88.78 ;
    RECT 65.525 88.02 65.745 88.78 ;
    RECT 66.225 88.02 66.445 88.78 ;
    RECT 66.925 88.02 67.14 88.78 ;
    RECT 67.62 88.02 67.84 88.78 ;
    RECT 68.32 88.02 69.235 88.78 ;
    RECT 69.715 88.02 69.935 88.78 ;
    RECT 70.415 88.02 70.635 88.78 ;
    RECT 71.115 88.02 71.335 88.78 ;
    RECT 71.815 88.02 72.035 88.78 ;
    RECT 72.515 88.02 72.735 88.78 ;
    RECT 73.215 88.02 73.435 88.78 ;
    RECT 73.915 88.02 74.835 88.78 ;
    RECT 75.315 88.02 75.535 88.78 ;
    RECT 76.015 88.02 76.225 88.78 ;
    RECT 76.705 88.02 76.92 88.78 ;
    RECT 77.4 88.02 77.62 88.78 ;
    RECT 78.1 88.02 78.32 88.78 ;
    RECT 78.8 88.02 79.02 88.78 ;
    RECT 79.5 88.02 81.115 88.78 ;
    RECT 81.595 88.02 81.815 88.78 ;
    RECT 82.295 88.02 82.515 88.78 ;
    RECT 82.995 88.02 83.055 88.78 ;
    RECT 83.055 87.93 83.335 88.87 ;
    RECT 83.335 88.02 83.505 88.78 ;
    RECT 26.71 87.26 26.88 88.02 ;
    RECT 26.88 87.17 27.16 88.11 ;
    RECT 27.16 87.26 27.32 88.02 ;
    RECT 27.8 87.26 28.02 88.02 ;
    RECT 28.5 87.26 28.72 88.02 ;
    RECT 29.2 87.26 30.815 88.02 ;
    RECT 31.295 87.26 31.515 88.02 ;
    RECT 31.995 87.26 32.21 88.02 ;
    RECT 32.69 87.26 32.91 88.02 ;
    RECT 33.39 87.26 33.61 88.02 ;
    RECT 34.09 87.26 34.31 88.02 ;
    RECT 34.79 87.26 35.005 88.02 ;
    RECT 35.485 87.26 36.405 88.02 ;
    RECT 36.885 87.26 37.105 88.02 ;
    RECT 37.585 87.26 37.8 88.02 ;
    RECT 38.28 87.26 38.5 88.02 ;
    RECT 38.98 87.26 39.2 88.02 ;
    RECT 39.68 87.26 39.895 88.02 ;
    RECT 40.375 87.26 40.595 88.02 ;
    RECT 41.075 87.26 41.995 88.02 ;
    RECT 42.475 87.26 42.69 88.02 ;
    RECT 43.17 87.26 43.39 88.02 ;
    RECT 43.87 87.26 44.09 88.02 ;
    RECT 44.57 87.26 44.79 88.02 ;
    RECT 45.27 87.26 45.485 88.02 ;
    RECT 45.965 87.26 46.185 88.02 ;
    RECT 46.665 87.26 47.58 88.02 ;
    RECT 48.06 87.26 48.28 88.02 ;
    RECT 48.76 87.26 48.98 88.02 ;
    RECT 49.46 87.26 49.68 88.02 ;
    RECT 50.16 87.26 50.375 88.02 ;
    RECT 50.855 87.26 51.775 88.02 ;
    RECT 52.255 87.26 53.17 88.02 ;
    RECT 53.65 87.26 53.87 88.02 ;
    RECT 54.35 87.26 54.57 88.02 ;
    RECT 55.05 87.26 55.265 88.02 ;
    RECT 55.745 87.26 55.965 88.02 ;
    RECT 56.445 87.26 56.665 88.02 ;
    RECT 57.145 87.26 58.06 88.02 ;
    RECT 58.54 87.26 59.46 88.02 ;
    RECT 59.94 87.26 60.16 88.02 ;
    RECT 60.64 87.26 60.855 88.02 ;
    RECT 61.335 87.26 61.555 88.02 ;
    RECT 62.035 87.26 62.25 88.02 ;
    RECT 62.73 87.26 63.65 88.02 ;
    RECT 64.13 87.26 64.345 88.02 ;
    RECT 64.825 87.26 65.045 88.02 ;
    RECT 65.525 87.26 65.745 88.02 ;
    RECT 66.225 87.26 66.445 88.02 ;
    RECT 66.925 87.26 67.14 88.02 ;
    RECT 67.62 87.26 67.84 88.02 ;
    RECT 68.32 87.26 69.235 88.02 ;
    RECT 69.715 87.26 69.935 88.02 ;
    RECT 70.415 87.26 70.635 88.02 ;
    RECT 71.115 87.26 71.335 88.02 ;
    RECT 71.815 87.26 72.035 88.02 ;
    RECT 72.515 87.26 72.735 88.02 ;
    RECT 73.215 87.26 73.435 88.02 ;
    RECT 73.915 87.26 74.835 88.02 ;
    RECT 75.315 87.26 75.535 88.02 ;
    RECT 76.015 87.26 76.225 88.02 ;
    RECT 76.705 87.26 76.92 88.02 ;
    RECT 77.4 87.26 77.62 88.02 ;
    RECT 78.1 87.26 78.32 88.02 ;
    RECT 78.8 87.26 79.02 88.02 ;
    RECT 79.5 87.26 81.115 88.02 ;
    RECT 81.595 87.26 81.815 88.02 ;
    RECT 82.295 87.26 82.515 88.02 ;
    RECT 82.995 87.26 83.055 88.02 ;
    RECT 83.055 87.17 83.335 88.11 ;
    RECT 83.335 87.26 83.505 88.02 ;
    RECT 26.71 109.3 26.88 110.77 ;
    RECT 26.88 109.205 27.16 110.77 ;
    RECT 27.16 109.3 27.32 110.77 ;
    RECT 27.8 109.3 28.02 110.77 ;
    RECT 28.5 109.3 28.72 110.77 ;
    RECT 29.2 109.3 30.815 110.77 ;
    RECT 31.295 109.3 31.515 110.77 ;
    RECT 31.995 109.3 32.21 110.77 ;
    RECT 32.69 109.3 32.91 110.77 ;
    RECT 33.39 109.3 33.61 110.77 ;
    RECT 34.09 109.3 34.31 110.77 ;
    RECT 34.79 109.3 35.005 110.77 ;
    RECT 35.485 109.3 36.405 110.77 ;
    RECT 36.885 109.3 37.105 110.77 ;
    RECT 37.585 109.3 37.8 110.77 ;
    RECT 38.28 109.3 38.5 110.77 ;
    RECT 38.98 109.3 39.2 110.77 ;
    RECT 39.68 109.3 39.895 110.77 ;
    RECT 40.375 109.3 40.595 110.77 ;
    RECT 41.075 109.3 41.995 110.77 ;
    RECT 42.475 109.3 42.69 110.77 ;
    RECT 43.17 109.3 43.39 110.77 ;
    RECT 43.87 109.3 44.09 110.77 ;
    RECT 44.57 109.3 44.79 110.77 ;
    RECT 45.27 109.3 45.485 110.77 ;
    RECT 45.965 109.3 46.185 110.77 ;
    RECT 46.665 109.3 47.58 110.77 ;
    RECT 48.06 109.3 48.28 110.77 ;
    RECT 48.76 109.3 48.98 110.77 ;
    RECT 49.46 109.3 49.68 110.77 ;
    RECT 50.16 109.3 50.375 110.77 ;
    RECT 50.855 109.3 51.775 110.77 ;
    RECT 52.255 109.3 53.17 110.77 ;
    RECT 53.65 109.3 53.87 110.77 ;
    RECT 54.35 109.3 54.57 110.77 ;
    RECT 55.05 109.3 55.265 110.77 ;
    RECT 55.745 109.3 55.965 110.77 ;
    RECT 56.445 109.3 56.665 110.77 ;
    RECT 57.145 109.3 58.06 110.77 ;
    RECT 58.54 109.3 59.46 110.77 ;
    RECT 59.94 109.3 60.16 110.77 ;
    RECT 60.64 109.3 60.855 110.77 ;
    RECT 61.335 109.3 61.555 110.77 ;
    RECT 62.035 109.3 62.25 110.77 ;
    RECT 62.73 109.3 63.65 110.77 ;
    RECT 64.13 109.3 64.345 110.77 ;
    RECT 64.825 109.3 65.045 110.77 ;
    RECT 65.525 109.3 65.745 110.77 ;
    RECT 66.225 109.3 66.445 110.77 ;
    RECT 66.925 109.3 67.14 110.77 ;
    RECT 67.62 109.3 67.84 110.77 ;
    RECT 68.32 109.3 69.235 110.77 ;
    RECT 69.715 109.3 69.935 110.77 ;
    RECT 70.415 109.3 70.635 110.77 ;
    RECT 71.115 109.3 71.335 110.77 ;
    RECT 71.815 109.3 72.035 110.77 ;
    RECT 72.515 109.3 72.735 110.77 ;
    RECT 73.215 109.3 73.435 110.77 ;
    RECT 73.915 109.3 74.835 110.77 ;
    RECT 75.315 109.3 75.535 110.77 ;
    RECT 76.015 109.3 76.225 110.77 ;
    RECT 76.705 109.3 76.92 110.77 ;
    RECT 77.4 109.3 77.62 110.77 ;
    RECT 78.1 109.3 78.32 110.77 ;
    RECT 78.8 109.3 79.02 110.77 ;
    RECT 79.5 109.3 81.115 110.77 ;
    RECT 81.595 109.3 81.815 110.77 ;
    RECT 82.295 109.3 82.515 110.77 ;
    RECT 82.995 109.3 83.505 110.77 ;
    RECT 26.71 108.54 26.88 109.3 ;
    RECT 26.88 108.45 27.16 109.39 ;
    RECT 27.16 108.54 27.32 109.3 ;
    RECT 27.8 108.54 28.02 109.3 ;
    RECT 28.5 108.54 28.72 109.3 ;
    RECT 29.2 108.54 30.815 109.3 ;
    RECT 31.295 108.54 31.515 109.3 ;
    RECT 31.995 108.54 32.21 109.3 ;
    RECT 32.69 108.54 32.91 109.3 ;
    RECT 33.39 108.54 33.61 109.3 ;
    RECT 34.09 108.54 34.31 109.3 ;
    RECT 34.79 108.54 35.005 109.3 ;
    RECT 35.485 108.54 36.405 109.3 ;
    RECT 36.885 108.54 37.105 109.3 ;
    RECT 37.585 108.54 37.8 109.3 ;
    RECT 38.28 108.54 38.5 109.3 ;
    RECT 38.98 108.54 39.2 109.3 ;
    RECT 39.68 108.54 39.895 109.3 ;
    RECT 40.375 108.54 40.595 109.3 ;
    RECT 41.075 108.54 41.995 109.3 ;
    RECT 42.475 108.54 42.69 109.3 ;
    RECT 43.17 108.54 43.39 109.3 ;
    RECT 43.87 108.54 44.09 109.3 ;
    RECT 44.57 108.54 44.79 109.3 ;
    RECT 45.27 108.54 45.485 109.3 ;
    RECT 45.965 108.54 46.185 109.3 ;
    RECT 46.665 108.54 47.58 109.3 ;
    RECT 48.06 108.54 48.28 109.3 ;
    RECT 48.76 108.54 48.98 109.3 ;
    RECT 49.46 108.54 49.68 109.3 ;
    RECT 50.16 108.54 50.375 109.3 ;
    RECT 50.855 108.54 51.775 109.3 ;
    RECT 52.255 108.54 53.17 109.3 ;
    RECT 53.65 108.54 53.87 109.3 ;
    RECT 54.35 108.54 54.57 109.3 ;
    RECT 55.05 108.54 55.265 109.3 ;
    RECT 55.745 108.54 55.965 109.3 ;
    RECT 56.445 108.54 56.665 109.3 ;
    RECT 57.145 108.54 58.06 109.3 ;
    RECT 58.54 108.54 59.46 109.3 ;
    RECT 59.94 108.54 60.16 109.3 ;
    RECT 60.64 108.54 60.855 109.3 ;
    RECT 61.335 108.54 61.555 109.3 ;
    RECT 62.035 108.54 62.25 109.3 ;
    RECT 62.73 108.54 63.65 109.3 ;
    RECT 64.13 108.54 64.345 109.3 ;
    RECT 64.825 108.54 65.045 109.3 ;
    RECT 65.525 108.54 65.745 109.3 ;
    RECT 66.225 108.54 66.445 109.3 ;
    RECT 66.925 108.54 67.14 109.3 ;
    RECT 67.62 108.54 67.84 109.3 ;
    RECT 68.32 108.54 69.235 109.3 ;
    RECT 69.715 108.54 69.935 109.3 ;
    RECT 70.415 108.54 70.635 109.3 ;
    RECT 71.115 108.54 71.335 109.3 ;
    RECT 71.815 108.54 72.035 109.3 ;
    RECT 72.515 108.54 72.735 109.3 ;
    RECT 73.215 108.54 73.435 109.3 ;
    RECT 73.915 108.54 74.835 109.3 ;
    RECT 75.315 108.54 75.535 109.3 ;
    RECT 76.015 108.54 76.225 109.3 ;
    RECT 76.705 108.54 76.92 109.3 ;
    RECT 77.4 108.54 77.62 109.3 ;
    RECT 78.1 108.54 78.32 109.3 ;
    RECT 78.8 108.54 79.02 109.3 ;
    RECT 79.5 108.54 81.115 109.3 ;
    RECT 81.595 108.54 81.815 109.3 ;
    RECT 82.295 108.54 82.515 109.3 ;
    RECT 82.995 108.54 83.055 109.3 ;
    RECT 83.055 108.45 83.335 109.39 ;
    RECT 83.335 108.54 83.505 109.3 ;
    RECT 26.71 86.5 26.88 87.26 ;
    RECT 26.88 86.41 27.16 87.35 ;
    RECT 27.16 86.5 27.32 87.26 ;
    RECT 27.8 86.5 28.02 87.26 ;
    RECT 28.5 86.5 28.72 87.26 ;
    RECT 29.2 86.5 30.815 87.26 ;
    RECT 31.295 86.5 31.515 87.26 ;
    RECT 31.995 86.5 32.21 87.26 ;
    RECT 32.69 86.5 32.91 87.26 ;
    RECT 33.39 86.5 33.61 87.26 ;
    RECT 34.09 86.5 34.31 87.26 ;
    RECT 34.79 86.5 35.005 87.26 ;
    RECT 35.485 86.5 36.405 87.26 ;
    RECT 36.885 86.5 37.105 87.26 ;
    RECT 37.585 86.5 37.8 87.26 ;
    RECT 38.28 86.5 38.5 87.26 ;
    RECT 38.98 86.5 39.2 87.26 ;
    RECT 39.68 86.5 39.895 87.26 ;
    RECT 40.375 86.5 40.595 87.26 ;
    RECT 41.075 86.5 41.995 87.26 ;
    RECT 42.475 86.5 42.69 87.26 ;
    RECT 43.17 86.5 43.39 87.26 ;
    RECT 43.87 86.5 44.09 87.26 ;
    RECT 44.57 86.5 44.79 87.26 ;
    RECT 45.27 86.5 45.485 87.26 ;
    RECT 45.965 86.5 46.185 87.26 ;
    RECT 46.665 86.5 47.58 87.26 ;
    RECT 48.06 86.5 48.28 87.26 ;
    RECT 48.76 86.5 48.98 87.26 ;
    RECT 49.46 86.5 49.68 87.26 ;
    RECT 50.16 86.5 50.375 87.26 ;
    RECT 50.855 86.5 51.775 87.26 ;
    RECT 52.255 86.5 53.17 87.26 ;
    RECT 53.65 86.5 53.87 87.26 ;
    RECT 54.35 86.5 54.57 87.26 ;
    RECT 55.05 86.5 55.265 87.26 ;
    RECT 55.745 86.5 55.965 87.26 ;
    RECT 56.445 86.5 56.665 87.26 ;
    RECT 57.145 86.5 58.06 87.26 ;
    RECT 58.54 86.5 59.46 87.26 ;
    RECT 59.94 86.5 60.16 87.26 ;
    RECT 60.64 86.5 60.855 87.26 ;
    RECT 61.335 86.5 61.555 87.26 ;
    RECT 62.035 86.5 62.25 87.26 ;
    RECT 62.73 86.5 63.65 87.26 ;
    RECT 64.13 86.5 64.345 87.26 ;
    RECT 64.825 86.5 65.045 87.26 ;
    RECT 65.525 86.5 65.745 87.26 ;
    RECT 66.225 86.5 66.445 87.26 ;
    RECT 66.925 86.5 67.14 87.26 ;
    RECT 67.62 86.5 67.84 87.26 ;
    RECT 68.32 86.5 69.235 87.26 ;
    RECT 69.715 86.5 69.935 87.26 ;
    RECT 70.415 86.5 70.635 87.26 ;
    RECT 71.115 86.5 71.335 87.26 ;
    RECT 71.815 86.5 72.035 87.26 ;
    RECT 72.515 86.5 72.735 87.26 ;
    RECT 73.215 86.5 73.435 87.26 ;
    RECT 73.915 86.5 74.835 87.26 ;
    RECT 75.315 86.5 75.535 87.26 ;
    RECT 76.015 86.5 76.225 87.26 ;
    RECT 76.705 86.5 76.92 87.26 ;
    RECT 77.4 86.5 77.62 87.26 ;
    RECT 78.1 86.5 78.32 87.26 ;
    RECT 78.8 86.5 79.02 87.26 ;
    RECT 79.5 86.5 81.115 87.26 ;
    RECT 81.595 86.5 81.815 87.26 ;
    RECT 82.295 86.5 82.515 87.26 ;
    RECT 82.995 86.5 83.055 87.26 ;
    RECT 83.055 86.41 83.335 87.35 ;
    RECT 83.335 86.5 83.505 87.26 ;
    RECT 26.71 85.74 26.88 86.5 ;
    RECT 26.88 85.65 27.16 86.59 ;
    RECT 27.16 85.74 27.32 86.5 ;
    RECT 27.8 85.74 28.02 86.5 ;
    RECT 28.5 85.74 28.72 86.5 ;
    RECT 29.2 85.74 30.815 86.5 ;
    RECT 31.295 85.74 31.515 86.5 ;
    RECT 31.995 85.74 32.21 86.5 ;
    RECT 32.69 85.74 32.91 86.5 ;
    RECT 33.39 85.74 33.61 86.5 ;
    RECT 34.09 85.74 34.31 86.5 ;
    RECT 34.79 85.74 35.005 86.5 ;
    RECT 35.485 85.74 36.405 86.5 ;
    RECT 36.885 85.74 37.105 86.5 ;
    RECT 37.585 85.74 37.8 86.5 ;
    RECT 38.28 85.74 38.5 86.5 ;
    RECT 38.98 85.74 39.2 86.5 ;
    RECT 39.68 85.74 39.895 86.5 ;
    RECT 40.375 85.74 40.595 86.5 ;
    RECT 41.075 85.74 41.995 86.5 ;
    RECT 42.475 85.74 42.69 86.5 ;
    RECT 43.17 85.74 43.39 86.5 ;
    RECT 43.87 85.74 44.09 86.5 ;
    RECT 44.57 85.74 44.79 86.5 ;
    RECT 45.27 85.74 45.485 86.5 ;
    RECT 45.965 85.74 46.185 86.5 ;
    RECT 46.665 85.74 47.58 86.5 ;
    RECT 48.06 85.74 48.28 86.5 ;
    RECT 48.76 85.74 48.98 86.5 ;
    RECT 49.46 85.74 49.68 86.5 ;
    RECT 50.16 85.74 50.375 86.5 ;
    RECT 50.855 85.74 51.775 86.5 ;
    RECT 52.255 85.74 53.17 86.5 ;
    RECT 53.65 85.74 53.87 86.5 ;
    RECT 54.35 85.74 54.57 86.5 ;
    RECT 55.05 85.74 55.265 86.5 ;
    RECT 55.745 85.74 55.965 86.5 ;
    RECT 56.445 85.74 56.665 86.5 ;
    RECT 57.145 85.74 58.06 86.5 ;
    RECT 58.54 85.74 59.46 86.5 ;
    RECT 59.94 85.74 60.16 86.5 ;
    RECT 60.64 85.74 60.855 86.5 ;
    RECT 61.335 85.74 61.555 86.5 ;
    RECT 62.035 85.74 62.25 86.5 ;
    RECT 62.73 85.74 63.65 86.5 ;
    RECT 64.13 85.74 64.345 86.5 ;
    RECT 64.825 85.74 65.045 86.5 ;
    RECT 65.525 85.74 65.745 86.5 ;
    RECT 66.225 85.74 66.445 86.5 ;
    RECT 66.925 85.74 67.14 86.5 ;
    RECT 67.62 85.74 67.84 86.5 ;
    RECT 68.32 85.74 69.235 86.5 ;
    RECT 69.715 85.74 69.935 86.5 ;
    RECT 70.415 85.74 70.635 86.5 ;
    RECT 71.115 85.74 71.335 86.5 ;
    RECT 71.815 85.74 72.035 86.5 ;
    RECT 72.515 85.74 72.735 86.5 ;
    RECT 73.215 85.74 73.435 86.5 ;
    RECT 73.915 85.74 74.835 86.5 ;
    RECT 75.315 85.74 75.535 86.5 ;
    RECT 76.015 85.74 76.225 86.5 ;
    RECT 76.705 85.74 76.92 86.5 ;
    RECT 77.4 85.74 77.62 86.5 ;
    RECT 78.1 85.74 78.32 86.5 ;
    RECT 78.8 85.74 79.02 86.5 ;
    RECT 79.5 85.74 81.115 86.5 ;
    RECT 81.595 85.74 81.815 86.5 ;
    RECT 82.295 85.74 82.515 86.5 ;
    RECT 82.995 85.74 83.055 86.5 ;
    RECT 83.055 85.65 83.335 86.59 ;
    RECT 83.335 85.74 83.505 86.5 ;
    RECT 26.71 84.98 26.88 85.74 ;
    RECT 26.88 84.89 27.16 85.83 ;
    RECT 27.16 84.98 27.32 85.74 ;
    RECT 27.8 84.98 28.02 85.74 ;
    RECT 28.5 84.98 28.72 85.74 ;
    RECT 29.2 84.98 30.815 85.74 ;
    RECT 31.295 84.98 31.515 85.74 ;
    RECT 31.995 84.98 32.21 85.74 ;
    RECT 32.69 84.98 32.91 85.74 ;
    RECT 33.39 84.98 33.61 85.74 ;
    RECT 34.09 84.98 34.31 85.74 ;
    RECT 34.79 84.98 35.005 85.74 ;
    RECT 35.485 84.98 36.405 85.74 ;
    RECT 36.885 84.98 37.105 85.74 ;
    RECT 37.585 84.98 37.8 85.74 ;
    RECT 38.28 84.98 38.5 85.74 ;
    RECT 38.98 84.98 39.2 85.74 ;
    RECT 39.68 84.98 39.895 85.74 ;
    RECT 40.375 84.98 40.595 85.74 ;
    RECT 41.075 84.98 41.995 85.74 ;
    RECT 42.475 84.98 42.69 85.74 ;
    RECT 43.17 84.98 43.39 85.74 ;
    RECT 43.87 84.98 44.09 85.74 ;
    RECT 44.57 84.98 44.79 85.74 ;
    RECT 45.27 84.98 45.485 85.74 ;
    RECT 45.965 84.98 46.185 85.74 ;
    RECT 46.665 84.98 47.58 85.74 ;
    RECT 48.06 84.98 48.28 85.74 ;
    RECT 48.76 84.98 48.98 85.74 ;
    RECT 49.46 84.98 49.68 85.74 ;
    RECT 50.16 84.98 50.375 85.74 ;
    RECT 50.855 84.98 51.775 85.74 ;
    RECT 52.255 84.98 53.17 85.74 ;
    RECT 53.65 84.98 53.87 85.74 ;
    RECT 54.35 84.98 54.57 85.74 ;
    RECT 55.05 84.98 55.265 85.74 ;
    RECT 55.745 84.98 55.965 85.74 ;
    RECT 56.445 84.98 56.665 85.74 ;
    RECT 57.145 84.98 58.06 85.74 ;
    RECT 58.54 84.98 59.46 85.74 ;
    RECT 59.94 84.98 60.16 85.74 ;
    RECT 60.64 84.98 60.855 85.74 ;
    RECT 61.335 84.98 61.555 85.74 ;
    RECT 62.035 84.98 62.25 85.74 ;
    RECT 62.73 84.98 63.65 85.74 ;
    RECT 64.13 84.98 64.345 85.74 ;
    RECT 64.825 84.98 65.045 85.74 ;
    RECT 65.525 84.98 65.745 85.74 ;
    RECT 66.225 84.98 66.445 85.74 ;
    RECT 66.925 84.98 67.14 85.74 ;
    RECT 67.62 84.98 67.84 85.74 ;
    RECT 68.32 84.98 69.235 85.74 ;
    RECT 69.715 84.98 69.935 85.74 ;
    RECT 70.415 84.98 70.635 85.74 ;
    RECT 71.115 84.98 71.335 85.74 ;
    RECT 71.815 84.98 72.035 85.74 ;
    RECT 72.515 84.98 72.735 85.74 ;
    RECT 73.215 84.98 73.435 85.74 ;
    RECT 73.915 84.98 74.835 85.74 ;
    RECT 75.315 84.98 75.535 85.74 ;
    RECT 76.015 84.98 76.225 85.74 ;
    RECT 76.705 84.98 76.92 85.74 ;
    RECT 77.4 84.98 77.62 85.74 ;
    RECT 78.1 84.98 78.32 85.74 ;
    RECT 78.8 84.98 79.02 85.74 ;
    RECT 79.5 84.98 81.115 85.74 ;
    RECT 81.595 84.98 81.815 85.74 ;
    RECT 82.295 84.98 82.515 85.74 ;
    RECT 82.995 84.98 83.055 85.74 ;
    RECT 83.055 84.89 83.335 85.83 ;
    RECT 83.335 84.98 83.505 85.74 ;
    RECT 26.71 84.22 26.88 84.98 ;
    RECT 26.88 84.13 27.16 85.07 ;
    RECT 27.16 84.22 27.32 84.98 ;
    RECT 27.8 84.22 28.02 84.98 ;
    RECT 28.5 84.22 28.72 84.98 ;
    RECT 29.2 84.22 30.815 84.98 ;
    RECT 31.295 84.22 31.515 84.98 ;
    RECT 31.995 84.22 32.21 84.98 ;
    RECT 32.69 84.22 32.91 84.98 ;
    RECT 33.39 84.22 33.61 84.98 ;
    RECT 34.09 84.22 34.31 84.98 ;
    RECT 34.79 84.22 35.005 84.98 ;
    RECT 35.485 84.22 36.405 84.98 ;
    RECT 36.885 84.22 37.105 84.98 ;
    RECT 37.585 84.22 37.8 84.98 ;
    RECT 38.28 84.22 38.5 84.98 ;
    RECT 38.98 84.22 39.2 84.98 ;
    RECT 39.68 84.22 39.895 84.98 ;
    RECT 40.375 84.22 40.595 84.98 ;
    RECT 41.075 84.22 41.995 84.98 ;
    RECT 42.475 84.22 42.69 84.98 ;
    RECT 43.17 84.22 43.39 84.98 ;
    RECT 43.87 84.22 44.09 84.98 ;
    RECT 44.57 84.22 44.79 84.98 ;
    RECT 45.27 84.22 45.485 84.98 ;
    RECT 45.965 84.22 46.185 84.98 ;
    RECT 46.665 84.22 47.58 84.98 ;
    RECT 48.06 84.22 48.28 84.98 ;
    RECT 48.76 84.22 48.98 84.98 ;
    RECT 49.46 84.22 49.68 84.98 ;
    RECT 50.16 84.22 50.375 84.98 ;
    RECT 50.855 84.22 51.775 84.98 ;
    RECT 52.255 84.22 53.17 84.98 ;
    RECT 53.65 84.22 53.87 84.98 ;
    RECT 54.35 84.22 54.57 84.98 ;
    RECT 55.05 84.22 55.265 84.98 ;
    RECT 55.745 84.22 55.965 84.98 ;
    RECT 56.445 84.22 56.665 84.98 ;
    RECT 57.145 84.22 58.06 84.98 ;
    RECT 58.54 84.22 59.46 84.98 ;
    RECT 59.94 84.22 60.16 84.98 ;
    RECT 60.64 84.22 60.855 84.98 ;
    RECT 61.335 84.22 61.555 84.98 ;
    RECT 62.035 84.22 62.25 84.98 ;
    RECT 62.73 84.22 63.65 84.98 ;
    RECT 64.13 84.22 64.345 84.98 ;
    RECT 64.825 84.22 65.045 84.98 ;
    RECT 65.525 84.22 65.745 84.98 ;
    RECT 66.225 84.22 66.445 84.98 ;
    RECT 66.925 84.22 67.14 84.98 ;
    RECT 67.62 84.22 67.84 84.98 ;
    RECT 68.32 84.22 69.235 84.98 ;
    RECT 69.715 84.22 69.935 84.98 ;
    RECT 70.415 84.22 70.635 84.98 ;
    RECT 71.115 84.22 71.335 84.98 ;
    RECT 71.815 84.22 72.035 84.98 ;
    RECT 72.515 84.22 72.735 84.98 ;
    RECT 73.215 84.22 73.435 84.98 ;
    RECT 73.915 84.22 74.835 84.98 ;
    RECT 75.315 84.22 75.535 84.98 ;
    RECT 76.015 84.22 76.225 84.98 ;
    RECT 76.705 84.22 76.92 84.98 ;
    RECT 77.4 84.22 77.62 84.98 ;
    RECT 78.1 84.22 78.32 84.98 ;
    RECT 78.8 84.22 79.02 84.98 ;
    RECT 79.5 84.22 81.115 84.98 ;
    RECT 81.595 84.22 81.815 84.98 ;
    RECT 82.295 84.22 82.515 84.98 ;
    RECT 82.995 84.22 83.055 84.98 ;
    RECT 83.055 84.13 83.335 85.07 ;
    RECT 83.335 84.22 83.505 84.98 ;
    RECT 26.71 83.46 26.88 84.22 ;
    RECT 26.88 83.37 27.16 84.31 ;
    RECT 27.16 83.46 27.32 84.22 ;
    RECT 27.8 83.46 28.02 84.22 ;
    RECT 28.5 83.46 28.72 84.22 ;
    RECT 29.2 83.46 30.815 84.22 ;
    RECT 31.295 83.46 31.515 84.22 ;
    RECT 31.995 83.46 32.21 84.22 ;
    RECT 32.69 83.46 32.91 84.22 ;
    RECT 33.39 83.46 33.61 84.22 ;
    RECT 34.09 83.46 34.31 84.22 ;
    RECT 34.79 83.46 35.005 84.22 ;
    RECT 35.485 83.46 36.405 84.22 ;
    RECT 36.885 83.46 37.105 84.22 ;
    RECT 37.585 83.46 37.8 84.22 ;
    RECT 38.28 83.46 38.5 84.22 ;
    RECT 38.98 83.46 39.2 84.22 ;
    RECT 39.68 83.46 39.895 84.22 ;
    RECT 40.375 83.46 40.595 84.22 ;
    RECT 41.075 83.46 41.995 84.22 ;
    RECT 42.475 83.46 42.69 84.22 ;
    RECT 43.17 83.46 43.39 84.22 ;
    RECT 43.87 83.46 44.09 84.22 ;
    RECT 44.57 83.46 44.79 84.22 ;
    RECT 45.27 83.46 45.485 84.22 ;
    RECT 45.965 83.46 46.185 84.22 ;
    RECT 46.665 83.46 47.58 84.22 ;
    RECT 48.06 83.46 48.28 84.22 ;
    RECT 48.76 83.46 48.98 84.22 ;
    RECT 49.46 83.46 49.68 84.22 ;
    RECT 50.16 83.46 50.375 84.22 ;
    RECT 50.855 83.46 51.775 84.22 ;
    RECT 52.255 83.46 53.17 84.22 ;
    RECT 53.65 83.46 53.87 84.22 ;
    RECT 54.35 83.46 54.57 84.22 ;
    RECT 55.05 83.46 55.265 84.22 ;
    RECT 55.745 83.46 55.965 84.22 ;
    RECT 56.445 83.46 56.665 84.22 ;
    RECT 57.145 83.46 58.06 84.22 ;
    RECT 58.54 83.46 59.46 84.22 ;
    RECT 59.94 83.46 60.16 84.22 ;
    RECT 60.64 83.46 60.855 84.22 ;
    RECT 61.335 83.46 61.555 84.22 ;
    RECT 62.035 83.46 62.25 84.22 ;
    RECT 62.73 83.46 63.65 84.22 ;
    RECT 64.13 83.46 64.345 84.22 ;
    RECT 64.825 83.46 65.045 84.22 ;
    RECT 65.525 83.46 65.745 84.22 ;
    RECT 66.225 83.46 66.445 84.22 ;
    RECT 66.925 83.46 67.14 84.22 ;
    RECT 67.62 83.46 67.84 84.22 ;
    RECT 68.32 83.46 69.235 84.22 ;
    RECT 69.715 83.46 69.935 84.22 ;
    RECT 70.415 83.46 70.635 84.22 ;
    RECT 71.115 83.46 71.335 84.22 ;
    RECT 71.815 83.46 72.035 84.22 ;
    RECT 72.515 83.46 72.735 84.22 ;
    RECT 73.215 83.46 73.435 84.22 ;
    RECT 73.915 83.46 74.835 84.22 ;
    RECT 75.315 83.46 75.535 84.22 ;
    RECT 76.015 83.46 76.225 84.22 ;
    RECT 76.705 83.46 76.92 84.22 ;
    RECT 77.4 83.46 77.62 84.22 ;
    RECT 78.1 83.46 78.32 84.22 ;
    RECT 78.8 83.46 79.02 84.22 ;
    RECT 79.5 83.46 81.115 84.22 ;
    RECT 81.595 83.46 81.815 84.22 ;
    RECT 82.295 83.46 82.515 84.22 ;
    RECT 82.995 83.46 83.055 84.22 ;
    RECT 83.055 83.37 83.335 84.31 ;
    RECT 83.335 83.46 83.505 84.22 ;
    RECT 26.71 82.7 26.88 83.46 ;
    RECT 26.88 82.61 27.16 83.55 ;
    RECT 27.16 82.7 27.32 83.46 ;
    RECT 27.8 82.7 28.02 83.46 ;
    RECT 28.5 82.7 28.72 83.46 ;
    RECT 29.2 82.7 30.815 83.46 ;
    RECT 31.295 82.7 31.515 83.46 ;
    RECT 31.995 82.7 32.21 83.46 ;
    RECT 32.69 82.7 32.91 83.46 ;
    RECT 33.39 82.7 33.61 83.46 ;
    RECT 34.09 82.7 34.31 83.46 ;
    RECT 34.79 82.7 35.005 83.46 ;
    RECT 35.485 82.7 36.405 83.46 ;
    RECT 36.885 82.7 37.105 83.46 ;
    RECT 37.585 82.7 37.8 83.46 ;
    RECT 38.28 82.7 38.5 83.46 ;
    RECT 38.98 82.7 39.2 83.46 ;
    RECT 39.68 82.7 39.895 83.46 ;
    RECT 40.375 82.7 40.595 83.46 ;
    RECT 41.075 82.7 41.995 83.46 ;
    RECT 42.475 82.7 42.69 83.46 ;
    RECT 43.17 82.7 43.39 83.46 ;
    RECT 43.87 82.7 44.09 83.46 ;
    RECT 44.57 82.7 44.79 83.46 ;
    RECT 45.27 82.7 45.485 83.46 ;
    RECT 45.965 82.7 46.185 83.46 ;
    RECT 46.665 82.7 47.58 83.46 ;
    RECT 48.06 82.7 48.28 83.46 ;
    RECT 48.76 82.7 48.98 83.46 ;
    RECT 49.46 82.7 49.68 83.46 ;
    RECT 50.16 82.7 50.375 83.46 ;
    RECT 50.855 82.7 51.775 83.46 ;
    RECT 52.255 82.7 53.17 83.46 ;
    RECT 53.65 82.7 53.87 83.46 ;
    RECT 54.35 82.7 54.57 83.46 ;
    RECT 55.05 82.7 55.265 83.46 ;
    RECT 55.745 82.7 55.965 83.46 ;
    RECT 56.445 82.7 56.665 83.46 ;
    RECT 57.145 82.7 58.06 83.46 ;
    RECT 58.54 82.7 59.46 83.46 ;
    RECT 59.94 82.7 60.16 83.46 ;
    RECT 60.64 82.7 60.855 83.46 ;
    RECT 61.335 82.7 61.555 83.46 ;
    RECT 62.035 82.7 62.25 83.46 ;
    RECT 62.73 82.7 63.65 83.46 ;
    RECT 64.13 82.7 64.345 83.46 ;
    RECT 64.825 82.7 65.045 83.46 ;
    RECT 65.525 82.7 65.745 83.46 ;
    RECT 66.225 82.7 66.445 83.46 ;
    RECT 66.925 82.7 67.14 83.46 ;
    RECT 67.62 82.7 67.84 83.46 ;
    RECT 68.32 82.7 69.235 83.46 ;
    RECT 69.715 82.7 69.935 83.46 ;
    RECT 70.415 82.7 70.635 83.46 ;
    RECT 71.115 82.7 71.335 83.46 ;
    RECT 71.815 82.7 72.035 83.46 ;
    RECT 72.515 82.7 72.735 83.46 ;
    RECT 73.215 82.7 73.435 83.46 ;
    RECT 73.915 82.7 74.835 83.46 ;
    RECT 75.315 82.7 75.535 83.46 ;
    RECT 76.015 82.7 76.225 83.46 ;
    RECT 76.705 82.7 76.92 83.46 ;
    RECT 77.4 82.7 77.62 83.46 ;
    RECT 78.1 82.7 78.32 83.46 ;
    RECT 78.8 82.7 79.02 83.46 ;
    RECT 79.5 82.7 81.115 83.46 ;
    RECT 81.595 82.7 81.815 83.46 ;
    RECT 82.295 82.7 82.515 83.46 ;
    RECT 82.995 82.7 83.055 83.46 ;
    RECT 83.055 82.61 83.335 83.55 ;
    RECT 83.335 82.7 83.505 83.46 ;
    RECT 26.71 81.94 26.88 82.7 ;
    RECT 26.88 81.85 27.16 82.79 ;
    RECT 27.16 81.94 27.32 82.7 ;
    RECT 27.8 81.94 28.02 82.7 ;
    RECT 28.5 81.94 28.72 82.7 ;
    RECT 29.2 81.94 30.815 82.7 ;
    RECT 31.295 81.94 31.515 82.7 ;
    RECT 31.995 81.94 32.21 82.7 ;
    RECT 32.69 81.94 32.91 82.7 ;
    RECT 33.39 81.94 33.61 82.7 ;
    RECT 34.09 81.94 34.31 82.7 ;
    RECT 34.79 81.94 35.005 82.7 ;
    RECT 35.485 81.94 36.405 82.7 ;
    RECT 36.885 81.94 37.105 82.7 ;
    RECT 37.585 81.94 37.8 82.7 ;
    RECT 38.28 81.94 38.5 82.7 ;
    RECT 38.98 81.94 39.2 82.7 ;
    RECT 39.68 81.94 39.895 82.7 ;
    RECT 40.375 81.94 40.595 82.7 ;
    RECT 41.075 81.94 41.995 82.7 ;
    RECT 42.475 81.94 42.69 82.7 ;
    RECT 43.17 81.94 43.39 82.7 ;
    RECT 43.87 81.94 44.09 82.7 ;
    RECT 44.57 81.94 44.79 82.7 ;
    RECT 45.27 81.94 45.485 82.7 ;
    RECT 45.965 81.94 46.185 82.7 ;
    RECT 46.665 81.94 47.58 82.7 ;
    RECT 48.06 81.94 48.28 82.7 ;
    RECT 48.76 81.94 48.98 82.7 ;
    RECT 49.46 81.94 49.68 82.7 ;
    RECT 50.16 81.94 50.375 82.7 ;
    RECT 50.855 81.94 51.775 82.7 ;
    RECT 52.255 81.94 53.17 82.7 ;
    RECT 53.65 81.94 53.87 82.7 ;
    RECT 54.35 81.94 54.57 82.7 ;
    RECT 55.05 81.94 55.265 82.7 ;
    RECT 55.745 81.94 55.965 82.7 ;
    RECT 56.445 81.94 56.665 82.7 ;
    RECT 57.145 81.94 58.06 82.7 ;
    RECT 58.54 81.94 59.46 82.7 ;
    RECT 59.94 81.94 60.16 82.7 ;
    RECT 60.64 81.94 60.855 82.7 ;
    RECT 61.335 81.94 61.555 82.7 ;
    RECT 62.035 81.94 62.25 82.7 ;
    RECT 62.73 81.94 63.65 82.7 ;
    RECT 64.13 81.94 64.345 82.7 ;
    RECT 64.825 81.94 65.045 82.7 ;
    RECT 65.525 81.94 65.745 82.7 ;
    RECT 66.225 81.94 66.445 82.7 ;
    RECT 66.925 81.94 67.14 82.7 ;
    RECT 67.62 81.94 67.84 82.7 ;
    RECT 68.32 81.94 69.235 82.7 ;
    RECT 69.715 81.94 69.935 82.7 ;
    RECT 70.415 81.94 70.635 82.7 ;
    RECT 71.115 81.94 71.335 82.7 ;
    RECT 71.815 81.94 72.035 82.7 ;
    RECT 72.515 81.94 72.735 82.7 ;
    RECT 73.215 81.94 73.435 82.7 ;
    RECT 73.915 81.94 74.835 82.7 ;
    RECT 75.315 81.94 75.535 82.7 ;
    RECT 76.015 81.94 76.225 82.7 ;
    RECT 76.705 81.94 76.92 82.7 ;
    RECT 77.4 81.94 77.62 82.7 ;
    RECT 78.1 81.94 78.32 82.7 ;
    RECT 78.8 81.94 79.02 82.7 ;
    RECT 79.5 81.94 81.115 82.7 ;
    RECT 81.595 81.94 81.815 82.7 ;
    RECT 82.295 81.94 82.515 82.7 ;
    RECT 82.995 81.94 83.055 82.7 ;
    RECT 83.055 81.85 83.335 82.79 ;
    RECT 83.335 81.94 83.505 82.7 ;
    RECT 26.71 81.18 26.88 81.94 ;
    RECT 26.88 81.09 27.16 82.03 ;
    RECT 27.16 81.18 27.32 81.94 ;
    RECT 27.8 81.18 28.02 81.94 ;
    RECT 28.5 81.18 28.72 81.94 ;
    RECT 29.2 81.18 30.815 81.94 ;
    RECT 31.295 81.18 31.515 81.94 ;
    RECT 31.995 81.18 32.21 81.94 ;
    RECT 32.69 81.18 32.91 81.94 ;
    RECT 33.39 81.18 33.61 81.94 ;
    RECT 34.09 81.18 34.31 81.94 ;
    RECT 34.79 81.18 35.005 81.94 ;
    RECT 35.485 81.18 36.405 81.94 ;
    RECT 36.885 81.18 37.105 81.94 ;
    RECT 37.585 81.18 37.8 81.94 ;
    RECT 38.28 81.18 38.5 81.94 ;
    RECT 38.98 81.18 39.2 81.94 ;
    RECT 39.68 81.18 39.895 81.94 ;
    RECT 40.375 81.18 40.595 81.94 ;
    RECT 41.075 81.18 41.995 81.94 ;
    RECT 42.475 81.18 42.69 81.94 ;
    RECT 43.17 81.18 43.39 81.94 ;
    RECT 43.87 81.18 44.09 81.94 ;
    RECT 44.57 81.18 44.79 81.94 ;
    RECT 45.27 81.18 45.485 81.94 ;
    RECT 45.965 81.18 46.185 81.94 ;
    RECT 46.665 81.18 47.58 81.94 ;
    RECT 48.06 81.18 48.28 81.94 ;
    RECT 48.76 81.18 48.98 81.94 ;
    RECT 49.46 81.18 49.68 81.94 ;
    RECT 50.16 81.18 50.375 81.94 ;
    RECT 50.855 81.18 51.775 81.94 ;
    RECT 52.255 81.18 53.17 81.94 ;
    RECT 53.65 81.18 53.87 81.94 ;
    RECT 54.35 81.18 54.57 81.94 ;
    RECT 55.05 81.18 55.265 81.94 ;
    RECT 55.745 81.18 55.965 81.94 ;
    RECT 56.445 81.18 56.665 81.94 ;
    RECT 57.145 81.18 58.06 81.94 ;
    RECT 58.54 81.18 59.46 81.94 ;
    RECT 59.94 81.18 60.16 81.94 ;
    RECT 60.64 81.18 60.855 81.94 ;
    RECT 61.335 81.18 61.555 81.94 ;
    RECT 62.035 81.18 62.25 81.94 ;
    RECT 62.73 81.18 63.65 81.94 ;
    RECT 64.13 81.18 64.345 81.94 ;
    RECT 64.825 81.18 65.045 81.94 ;
    RECT 65.525 81.18 65.745 81.94 ;
    RECT 66.225 81.18 66.445 81.94 ;
    RECT 66.925 81.18 67.14 81.94 ;
    RECT 67.62 81.18 67.84 81.94 ;
    RECT 68.32 81.18 69.235 81.94 ;
    RECT 69.715 81.18 69.935 81.94 ;
    RECT 70.415 81.18 70.635 81.94 ;
    RECT 71.115 81.18 71.335 81.94 ;
    RECT 71.815 81.18 72.035 81.94 ;
    RECT 72.515 81.18 72.735 81.94 ;
    RECT 73.215 81.18 73.435 81.94 ;
    RECT 73.915 81.18 74.835 81.94 ;
    RECT 75.315 81.18 75.535 81.94 ;
    RECT 76.015 81.18 76.225 81.94 ;
    RECT 76.705 81.18 76.92 81.94 ;
    RECT 77.4 81.18 77.62 81.94 ;
    RECT 78.1 81.18 78.32 81.94 ;
    RECT 78.8 81.18 79.02 81.94 ;
    RECT 79.5 81.18 81.115 81.94 ;
    RECT 81.595 81.18 81.815 81.94 ;
    RECT 82.295 81.18 82.515 81.94 ;
    RECT 82.995 81.18 83.055 81.94 ;
    RECT 83.055 81.09 83.335 82.03 ;
    RECT 83.335 81.18 83.505 81.94 ;
    RECT 26.71 80.42 26.88 81.18 ;
    RECT 26.88 80.33 27.16 81.27 ;
    RECT 27.16 80.42 27.32 81.18 ;
    RECT 27.8 80.42 28.02 81.18 ;
    RECT 28.5 80.42 28.72 81.18 ;
    RECT 29.2 80.42 30.815 81.18 ;
    RECT 31.295 80.42 31.515 81.18 ;
    RECT 31.995 80.42 32.21 81.18 ;
    RECT 32.69 80.42 32.91 81.18 ;
    RECT 33.39 80.42 33.61 81.18 ;
    RECT 34.09 80.42 34.31 81.18 ;
    RECT 34.79 80.42 35.005 81.18 ;
    RECT 35.485 80.42 36.405 81.18 ;
    RECT 36.885 80.42 37.105 81.18 ;
    RECT 37.585 80.42 37.8 81.18 ;
    RECT 38.28 80.42 38.5 81.18 ;
    RECT 38.98 80.42 39.2 81.18 ;
    RECT 39.68 80.42 39.895 81.18 ;
    RECT 40.375 80.42 40.595 81.18 ;
    RECT 41.075 80.42 41.995 81.18 ;
    RECT 42.475 80.42 42.69 81.18 ;
    RECT 43.17 80.42 43.39 81.18 ;
    RECT 43.87 80.42 44.09 81.18 ;
    RECT 44.57 80.42 44.79 81.18 ;
    RECT 45.27 80.42 45.485 81.18 ;
    RECT 45.965 80.42 46.185 81.18 ;
    RECT 46.665 80.42 47.58 81.18 ;
    RECT 48.06 80.42 48.28 81.18 ;
    RECT 48.76 80.42 48.98 81.18 ;
    RECT 49.46 80.42 49.68 81.18 ;
    RECT 50.16 80.42 50.375 81.18 ;
    RECT 50.855 80.42 51.775 81.18 ;
    RECT 52.255 80.42 53.17 81.18 ;
    RECT 53.65 80.42 53.87 81.18 ;
    RECT 54.35 80.42 54.57 81.18 ;
    RECT 55.05 80.42 55.265 81.18 ;
    RECT 55.745 80.42 55.965 81.18 ;
    RECT 56.445 80.42 56.665 81.18 ;
    RECT 57.145 80.42 58.06 81.18 ;
    RECT 58.54 80.42 59.46 81.18 ;
    RECT 59.94 80.42 60.16 81.18 ;
    RECT 60.64 80.42 60.855 81.18 ;
    RECT 61.335 80.42 61.555 81.18 ;
    RECT 62.035 80.42 62.25 81.18 ;
    RECT 62.73 80.42 63.65 81.18 ;
    RECT 64.13 80.42 64.345 81.18 ;
    RECT 64.825 80.42 65.045 81.18 ;
    RECT 65.525 80.42 65.745 81.18 ;
    RECT 66.225 80.42 66.445 81.18 ;
    RECT 66.925 80.42 67.14 81.18 ;
    RECT 67.62 80.42 67.84 81.18 ;
    RECT 68.32 80.42 69.235 81.18 ;
    RECT 69.715 80.42 69.935 81.18 ;
    RECT 70.415 80.42 70.635 81.18 ;
    RECT 71.115 80.42 71.335 81.18 ;
    RECT 71.815 80.42 72.035 81.18 ;
    RECT 72.515 80.42 72.735 81.18 ;
    RECT 73.215 80.42 73.435 81.18 ;
    RECT 73.915 80.42 74.835 81.18 ;
    RECT 75.315 80.42 75.535 81.18 ;
    RECT 76.015 80.42 76.225 81.18 ;
    RECT 76.705 80.42 76.92 81.18 ;
    RECT 77.4 80.42 77.62 81.18 ;
    RECT 78.1 80.42 78.32 81.18 ;
    RECT 78.8 80.42 79.02 81.18 ;
    RECT 79.5 80.42 81.115 81.18 ;
    RECT 81.595 80.42 81.815 81.18 ;
    RECT 82.295 80.42 82.515 81.18 ;
    RECT 82.995 80.42 83.055 81.18 ;
    RECT 83.055 80.33 83.335 81.27 ;
    RECT 83.335 80.42 83.505 81.18 ;
    RECT 26.71 79.66 26.88 80.42 ;
    RECT 26.88 79.57 27.16 80.51 ;
    RECT 27.16 79.66 27.32 80.42 ;
    RECT 27.8 79.66 28.02 80.42 ;
    RECT 28.5 79.66 28.72 80.42 ;
    RECT 29.2 79.66 30.815 80.42 ;
    RECT 31.295 79.66 31.515 80.42 ;
    RECT 31.995 79.66 32.21 80.42 ;
    RECT 32.69 79.66 32.91 80.42 ;
    RECT 33.39 79.66 33.61 80.42 ;
    RECT 34.09 79.66 34.31 80.42 ;
    RECT 34.79 79.66 35.005 80.42 ;
    RECT 35.485 79.66 36.405 80.42 ;
    RECT 36.885 79.66 37.105 80.42 ;
    RECT 37.585 79.66 37.8 80.42 ;
    RECT 38.28 79.66 38.5 80.42 ;
    RECT 38.98 79.66 39.2 80.42 ;
    RECT 39.68 79.66 39.895 80.42 ;
    RECT 40.375 79.66 40.595 80.42 ;
    RECT 41.075 79.66 41.995 80.42 ;
    RECT 42.475 79.66 42.69 80.42 ;
    RECT 43.17 79.66 43.39 80.42 ;
    RECT 43.87 79.66 44.09 80.42 ;
    RECT 44.57 79.66 44.79 80.42 ;
    RECT 45.27 79.66 45.485 80.42 ;
    RECT 45.965 79.66 46.185 80.42 ;
    RECT 46.665 79.66 47.58 80.42 ;
    RECT 48.06 79.66 48.28 80.42 ;
    RECT 48.76 79.66 48.98 80.42 ;
    RECT 49.46 79.66 49.68 80.42 ;
    RECT 50.16 79.66 50.375 80.42 ;
    RECT 50.855 79.66 51.775 80.42 ;
    RECT 52.255 79.66 53.17 80.42 ;
    RECT 53.65 79.66 53.87 80.42 ;
    RECT 54.35 79.66 54.57 80.42 ;
    RECT 55.05 79.66 55.265 80.42 ;
    RECT 55.745 79.66 55.965 80.42 ;
    RECT 56.445 79.66 56.665 80.42 ;
    RECT 57.145 79.66 58.06 80.42 ;
    RECT 58.54 79.66 59.46 80.42 ;
    RECT 59.94 79.66 60.16 80.42 ;
    RECT 60.64 79.66 60.855 80.42 ;
    RECT 61.335 79.66 61.555 80.42 ;
    RECT 62.035 79.66 62.25 80.42 ;
    RECT 62.73 79.66 63.65 80.42 ;
    RECT 64.13 79.66 64.345 80.42 ;
    RECT 64.825 79.66 65.045 80.42 ;
    RECT 65.525 79.66 65.745 80.42 ;
    RECT 66.225 79.66 66.445 80.42 ;
    RECT 66.925 79.66 67.14 80.42 ;
    RECT 67.62 79.66 67.84 80.42 ;
    RECT 68.32 79.66 69.235 80.42 ;
    RECT 69.715 79.66 69.935 80.42 ;
    RECT 70.415 79.66 70.635 80.42 ;
    RECT 71.115 79.66 71.335 80.42 ;
    RECT 71.815 79.66 72.035 80.42 ;
    RECT 72.515 79.66 72.735 80.42 ;
    RECT 73.215 79.66 73.435 80.42 ;
    RECT 73.915 79.66 74.835 80.42 ;
    RECT 75.315 79.66 75.535 80.42 ;
    RECT 76.015 79.66 76.225 80.42 ;
    RECT 76.705 79.66 76.92 80.42 ;
    RECT 77.4 79.66 77.62 80.42 ;
    RECT 78.1 79.66 78.32 80.42 ;
    RECT 78.8 79.66 79.02 80.42 ;
    RECT 79.5 79.66 81.115 80.42 ;
    RECT 81.595 79.66 81.815 80.42 ;
    RECT 82.295 79.66 82.515 80.42 ;
    RECT 82.995 79.66 83.055 80.42 ;
    RECT 83.055 79.57 83.335 80.51 ;
    RECT 83.335 79.66 83.505 80.42 ;
    RECT 26.71 78.9 26.88 79.66 ;
    RECT 26.88 78.81 27.16 79.75 ;
    RECT 27.16 78.9 27.32 79.66 ;
    RECT 27.8 78.9 28.02 79.66 ;
    RECT 28.5 78.9 28.72 79.66 ;
    RECT 29.2 78.9 30.815 79.66 ;
    RECT 31.295 78.9 31.515 79.66 ;
    RECT 31.995 78.9 32.21 79.66 ;
    RECT 32.69 78.9 32.91 79.66 ;
    RECT 33.39 78.9 33.61 79.66 ;
    RECT 34.09 78.9 34.31 79.66 ;
    RECT 34.79 78.9 35.005 79.66 ;
    RECT 35.485 78.9 36.405 79.66 ;
    RECT 36.885 78.9 37.105 79.66 ;
    RECT 37.585 78.9 37.8 79.66 ;
    RECT 38.28 78.9 38.5 79.66 ;
    RECT 38.98 78.9 39.2 79.66 ;
    RECT 39.68 78.9 39.895 79.66 ;
    RECT 40.375 78.9 40.595 79.66 ;
    RECT 41.075 78.9 41.995 79.66 ;
    RECT 42.475 78.9 42.69 79.66 ;
    RECT 43.17 78.9 43.39 79.66 ;
    RECT 43.87 78.9 44.09 79.66 ;
    RECT 44.57 78.9 44.79 79.66 ;
    RECT 45.27 78.9 45.485 79.66 ;
    RECT 45.965 78.9 46.185 79.66 ;
    RECT 46.665 78.9 47.58 79.66 ;
    RECT 48.06 78.9 48.28 79.66 ;
    RECT 48.76 78.9 48.98 79.66 ;
    RECT 49.46 78.9 49.68 79.66 ;
    RECT 50.16 78.9 50.375 79.66 ;
    RECT 50.855 78.9 51.775 79.66 ;
    RECT 52.255 78.9 53.17 79.66 ;
    RECT 53.65 78.9 53.87 79.66 ;
    RECT 54.35 78.9 54.57 79.66 ;
    RECT 55.05 78.9 55.265 79.66 ;
    RECT 55.745 78.9 55.965 79.66 ;
    RECT 56.445 78.9 56.665 79.66 ;
    RECT 57.145 78.9 58.06 79.66 ;
    RECT 58.54 78.9 59.46 79.66 ;
    RECT 59.94 78.9 60.16 79.66 ;
    RECT 60.64 78.9 60.855 79.66 ;
    RECT 61.335 78.9 61.555 79.66 ;
    RECT 62.035 78.9 62.25 79.66 ;
    RECT 62.73 78.9 63.65 79.66 ;
    RECT 64.13 78.9 64.345 79.66 ;
    RECT 64.825 78.9 65.045 79.66 ;
    RECT 65.525 78.9 65.745 79.66 ;
    RECT 66.225 78.9 66.445 79.66 ;
    RECT 66.925 78.9 67.14 79.66 ;
    RECT 67.62 78.9 67.84 79.66 ;
    RECT 68.32 78.9 69.235 79.66 ;
    RECT 69.715 78.9 69.935 79.66 ;
    RECT 70.415 78.9 70.635 79.66 ;
    RECT 71.115 78.9 71.335 79.66 ;
    RECT 71.815 78.9 72.035 79.66 ;
    RECT 72.515 78.9 72.735 79.66 ;
    RECT 73.215 78.9 73.435 79.66 ;
    RECT 73.915 78.9 74.835 79.66 ;
    RECT 75.315 78.9 75.535 79.66 ;
    RECT 76.015 78.9 76.225 79.66 ;
    RECT 76.705 78.9 76.92 79.66 ;
    RECT 77.4 78.9 77.62 79.66 ;
    RECT 78.1 78.9 78.32 79.66 ;
    RECT 78.8 78.9 79.02 79.66 ;
    RECT 79.5 78.9 81.115 79.66 ;
    RECT 81.595 78.9 81.815 79.66 ;
    RECT 82.295 78.9 82.515 79.66 ;
    RECT 82.995 78.9 83.055 79.66 ;
    RECT 83.055 78.81 83.335 79.75 ;
    RECT 83.335 78.9 83.505 79.66 ;
    RECT 26.71 78.14 26.88 78.9 ;
    RECT 26.88 78.05 27.16 78.99 ;
    RECT 27.16 78.14 27.32 78.9 ;
    RECT 27.8 78.14 28.02 78.9 ;
    RECT 28.5 78.14 28.72 78.9 ;
    RECT 29.2 78.14 30.815 78.9 ;
    RECT 31.295 78.14 31.515 78.9 ;
    RECT 31.995 78.14 32.21 78.9 ;
    RECT 32.69 78.14 32.91 78.9 ;
    RECT 33.39 78.14 33.61 78.9 ;
    RECT 34.09 78.14 34.31 78.9 ;
    RECT 34.79 78.14 35.005 78.9 ;
    RECT 35.485 78.14 36.405 78.9 ;
    RECT 36.885 78.14 37.105 78.9 ;
    RECT 37.585 78.14 37.8 78.9 ;
    RECT 38.28 78.14 38.5 78.9 ;
    RECT 38.98 78.14 39.2 78.9 ;
    RECT 39.68 78.14 39.895 78.9 ;
    RECT 40.375 78.14 40.595 78.9 ;
    RECT 41.075 78.14 41.995 78.9 ;
    RECT 42.475 78.14 42.69 78.9 ;
    RECT 43.17 78.14 43.39 78.9 ;
    RECT 43.87 78.14 44.09 78.9 ;
    RECT 44.57 78.14 44.79 78.9 ;
    RECT 45.27 78.14 45.485 78.9 ;
    RECT 45.965 78.14 46.185 78.9 ;
    RECT 46.665 78.14 47.58 78.9 ;
    RECT 48.06 78.14 48.28 78.9 ;
    RECT 48.76 78.14 48.98 78.9 ;
    RECT 49.46 78.14 49.68 78.9 ;
    RECT 50.16 78.14 50.375 78.9 ;
    RECT 50.855 78.14 51.775 78.9 ;
    RECT 52.255 78.14 53.17 78.9 ;
    RECT 53.65 78.14 53.87 78.9 ;
    RECT 54.35 78.14 54.57 78.9 ;
    RECT 55.05 78.14 55.265 78.9 ;
    RECT 55.745 78.14 55.965 78.9 ;
    RECT 56.445 78.14 56.665 78.9 ;
    RECT 57.145 78.14 58.06 78.9 ;
    RECT 58.54 78.14 59.46 78.9 ;
    RECT 59.94 78.14 60.16 78.9 ;
    RECT 60.64 78.14 60.855 78.9 ;
    RECT 61.335 78.14 61.555 78.9 ;
    RECT 62.035 78.14 62.25 78.9 ;
    RECT 62.73 78.14 63.65 78.9 ;
    RECT 64.13 78.14 64.345 78.9 ;
    RECT 64.825 78.14 65.045 78.9 ;
    RECT 65.525 78.14 65.745 78.9 ;
    RECT 66.225 78.14 66.445 78.9 ;
    RECT 66.925 78.14 67.14 78.9 ;
    RECT 67.62 78.14 67.84 78.9 ;
    RECT 68.32 78.14 69.235 78.9 ;
    RECT 69.715 78.14 69.935 78.9 ;
    RECT 70.415 78.14 70.635 78.9 ;
    RECT 71.115 78.14 71.335 78.9 ;
    RECT 71.815 78.14 72.035 78.9 ;
    RECT 72.515 78.14 72.735 78.9 ;
    RECT 73.215 78.14 73.435 78.9 ;
    RECT 73.915 78.14 74.835 78.9 ;
    RECT 75.315 78.14 75.535 78.9 ;
    RECT 76.015 78.14 76.225 78.9 ;
    RECT 76.705 78.14 76.92 78.9 ;
    RECT 77.4 78.14 77.62 78.9 ;
    RECT 78.1 78.14 78.32 78.9 ;
    RECT 78.8 78.14 79.02 78.9 ;
    RECT 79.5 78.14 81.115 78.9 ;
    RECT 81.595 78.14 81.815 78.9 ;
    RECT 82.295 78.14 82.515 78.9 ;
    RECT 82.995 78.14 83.055 78.9 ;
    RECT 83.055 78.05 83.335 78.99 ;
    RECT 83.335 78.14 83.505 78.9 ;
    RECT 26.71 77.38 26.88 78.14 ;
    RECT 26.88 77.29 27.16 78.23 ;
    RECT 27.16 77.38 27.32 78.14 ;
    RECT 27.8 77.38 28.02 78.14 ;
    RECT 28.5 77.38 28.72 78.14 ;
    RECT 29.2 77.38 30.815 78.14 ;
    RECT 31.295 77.38 31.515 78.14 ;
    RECT 31.995 77.38 32.21 78.14 ;
    RECT 32.69 77.38 32.91 78.14 ;
    RECT 33.39 77.38 33.61 78.14 ;
    RECT 34.09 77.38 34.31 78.14 ;
    RECT 34.79 77.38 35.005 78.14 ;
    RECT 35.485 77.38 36.405 78.14 ;
    RECT 36.885 77.38 37.105 78.14 ;
    RECT 37.585 77.38 37.8 78.14 ;
    RECT 38.28 77.38 38.5 78.14 ;
    RECT 38.98 77.38 39.2 78.14 ;
    RECT 39.68 77.38 39.895 78.14 ;
    RECT 40.375 77.38 40.595 78.14 ;
    RECT 41.075 77.38 41.995 78.14 ;
    RECT 42.475 77.38 42.69 78.14 ;
    RECT 43.17 77.38 43.39 78.14 ;
    RECT 43.87 77.38 44.09 78.14 ;
    RECT 44.57 77.38 44.79 78.14 ;
    RECT 45.27 77.38 45.485 78.14 ;
    RECT 45.965 77.38 46.185 78.14 ;
    RECT 46.665 77.38 47.58 78.14 ;
    RECT 48.06 77.38 48.28 78.14 ;
    RECT 48.76 77.38 48.98 78.14 ;
    RECT 49.46 77.38 49.68 78.14 ;
    RECT 50.16 77.38 50.375 78.14 ;
    RECT 50.855 77.38 51.775 78.14 ;
    RECT 52.255 77.38 53.17 78.14 ;
    RECT 53.65 77.38 53.87 78.14 ;
    RECT 54.35 77.38 54.57 78.14 ;
    RECT 55.05 77.38 55.265 78.14 ;
    RECT 55.745 77.38 55.965 78.14 ;
    RECT 56.445 77.38 56.665 78.14 ;
    RECT 57.145 77.38 58.06 78.14 ;
    RECT 58.54 77.38 59.46 78.14 ;
    RECT 59.94 77.38 60.16 78.14 ;
    RECT 60.64 77.38 60.855 78.14 ;
    RECT 61.335 77.38 61.555 78.14 ;
    RECT 62.035 77.38 62.25 78.14 ;
    RECT 62.73 77.38 63.65 78.14 ;
    RECT 64.13 77.38 64.345 78.14 ;
    RECT 64.825 77.38 65.045 78.14 ;
    RECT 65.525 77.38 65.745 78.14 ;
    RECT 66.225 77.38 66.445 78.14 ;
    RECT 66.925 77.38 67.14 78.14 ;
    RECT 67.62 77.38 67.84 78.14 ;
    RECT 68.32 77.38 69.235 78.14 ;
    RECT 69.715 77.38 69.935 78.14 ;
    RECT 70.415 77.38 70.635 78.14 ;
    RECT 71.115 77.38 71.335 78.14 ;
    RECT 71.815 77.38 72.035 78.14 ;
    RECT 72.515 77.38 72.735 78.14 ;
    RECT 73.215 77.38 73.435 78.14 ;
    RECT 73.915 77.38 74.835 78.14 ;
    RECT 75.315 77.38 75.535 78.14 ;
    RECT 76.015 77.38 76.225 78.14 ;
    RECT 76.705 77.38 76.92 78.14 ;
    RECT 77.4 77.38 77.62 78.14 ;
    RECT 78.1 77.38 78.32 78.14 ;
    RECT 78.8 77.38 79.02 78.14 ;
    RECT 79.5 77.38 81.115 78.14 ;
    RECT 81.595 77.38 81.815 78.14 ;
    RECT 82.295 77.38 82.515 78.14 ;
    RECT 82.995 77.38 83.055 78.14 ;
    RECT 83.055 77.29 83.335 78.23 ;
    RECT 83.335 77.38 83.505 78.14 ;
    RECT 26.71 76.62 26.88 77.38 ;
    RECT 26.88 76.53 27.16 77.47 ;
    RECT 27.16 76.62 27.32 77.38 ;
    RECT 27.8 76.62 28.02 77.38 ;
    RECT 28.5 76.62 28.72 77.38 ;
    RECT 29.2 76.62 30.815 77.38 ;
    RECT 31.295 76.62 31.515 77.38 ;
    RECT 31.995 76.62 32.21 77.38 ;
    RECT 32.69 76.62 32.91 77.38 ;
    RECT 33.39 76.62 33.61 77.38 ;
    RECT 34.09 76.62 34.31 77.38 ;
    RECT 34.79 76.62 35.005 77.38 ;
    RECT 35.485 76.62 36.405 77.38 ;
    RECT 36.885 76.62 37.105 77.38 ;
    RECT 37.585 76.62 37.8 77.38 ;
    RECT 38.28 76.62 38.5 77.38 ;
    RECT 38.98 76.62 39.2 77.38 ;
    RECT 39.68 76.62 39.895 77.38 ;
    RECT 40.375 76.62 40.595 77.38 ;
    RECT 41.075 76.62 41.995 77.38 ;
    RECT 42.475 76.62 42.69 77.38 ;
    RECT 43.17 76.62 43.39 77.38 ;
    RECT 43.87 76.62 44.09 77.38 ;
    RECT 44.57 76.62 44.79 77.38 ;
    RECT 45.27 76.62 45.485 77.38 ;
    RECT 45.965 76.62 46.185 77.38 ;
    RECT 46.665 76.62 47.58 77.38 ;
    RECT 48.06 76.62 48.28 77.38 ;
    RECT 48.76 76.62 48.98 77.38 ;
    RECT 49.46 76.62 49.68 77.38 ;
    RECT 50.16 76.62 50.375 77.38 ;
    RECT 50.855 76.62 51.775 77.38 ;
    RECT 52.255 76.62 53.17 77.38 ;
    RECT 53.65 76.62 53.87 77.38 ;
    RECT 54.35 76.62 54.57 77.38 ;
    RECT 55.05 76.62 55.265 77.38 ;
    RECT 55.745 76.62 55.965 77.38 ;
    RECT 56.445 76.62 56.665 77.38 ;
    RECT 57.145 76.62 58.06 77.38 ;
    RECT 58.54 76.62 59.46 77.38 ;
    RECT 59.94 76.62 60.16 77.38 ;
    RECT 60.64 76.62 60.855 77.38 ;
    RECT 61.335 76.62 61.555 77.38 ;
    RECT 62.035 76.62 62.25 77.38 ;
    RECT 62.73 76.62 63.65 77.38 ;
    RECT 64.13 76.62 64.345 77.38 ;
    RECT 64.825 76.62 65.045 77.38 ;
    RECT 65.525 76.62 65.745 77.38 ;
    RECT 66.225 76.62 66.445 77.38 ;
    RECT 66.925 76.62 67.14 77.38 ;
    RECT 67.62 76.62 67.84 77.38 ;
    RECT 68.32 76.62 69.235 77.38 ;
    RECT 69.715 76.62 69.935 77.38 ;
    RECT 70.415 76.62 70.635 77.38 ;
    RECT 71.115 76.62 71.335 77.38 ;
    RECT 71.815 76.62 72.035 77.38 ;
    RECT 72.515 76.62 72.735 77.38 ;
    RECT 73.215 76.62 73.435 77.38 ;
    RECT 73.915 76.62 74.835 77.38 ;
    RECT 75.315 76.62 75.535 77.38 ;
    RECT 76.015 76.62 76.225 77.38 ;
    RECT 76.705 76.62 76.92 77.38 ;
    RECT 77.4 76.62 77.62 77.38 ;
    RECT 78.1 76.62 78.32 77.38 ;
    RECT 78.8 76.62 79.02 77.38 ;
    RECT 79.5 76.62 81.115 77.38 ;
    RECT 81.595 76.62 81.815 77.38 ;
    RECT 82.295 76.62 82.515 77.38 ;
    RECT 82.995 76.62 83.055 77.38 ;
    RECT 83.055 76.53 83.335 77.47 ;
    RECT 83.335 76.62 83.505 77.38 ;
    RECT 26.71 75.86 26.88 76.62 ;
    RECT 26.88 75.77 27.16 76.71 ;
    RECT 27.16 75.86 27.32 76.62 ;
    RECT 27.8 75.86 28.02 76.62 ;
    RECT 28.5 75.86 28.72 76.62 ;
    RECT 29.2 75.86 30.815 76.62 ;
    RECT 31.295 75.86 31.515 76.62 ;
    RECT 31.995 75.86 32.21 76.62 ;
    RECT 32.69 75.86 32.91 76.62 ;
    RECT 33.39 75.86 33.61 76.62 ;
    RECT 34.09 75.86 34.31 76.62 ;
    RECT 34.79 75.86 35.005 76.62 ;
    RECT 35.485 75.86 36.405 76.62 ;
    RECT 36.885 75.86 37.105 76.62 ;
    RECT 37.585 75.86 37.8 76.62 ;
    RECT 38.28 75.86 38.5 76.62 ;
    RECT 38.98 75.86 39.2 76.62 ;
    RECT 39.68 75.86 39.895 76.62 ;
    RECT 40.375 75.86 40.595 76.62 ;
    RECT 41.075 75.86 41.995 76.62 ;
    RECT 42.475 75.86 42.69 76.62 ;
    RECT 43.17 75.86 43.39 76.62 ;
    RECT 43.87 75.86 44.09 76.62 ;
    RECT 44.57 75.86 44.79 76.62 ;
    RECT 45.27 75.86 45.485 76.62 ;
    RECT 45.965 75.86 46.185 76.62 ;
    RECT 46.665 75.86 47.58 76.62 ;
    RECT 48.06 75.86 48.28 76.62 ;
    RECT 48.76 75.86 48.98 76.62 ;
    RECT 49.46 75.86 49.68 76.62 ;
    RECT 50.16 75.86 50.375 76.62 ;
    RECT 50.855 75.86 51.775 76.62 ;
    RECT 52.255 75.86 53.17 76.62 ;
    RECT 53.65 75.86 53.87 76.62 ;
    RECT 54.35 75.86 54.57 76.62 ;
    RECT 55.05 75.86 55.265 76.62 ;
    RECT 55.745 75.86 55.965 76.62 ;
    RECT 56.445 75.86 56.665 76.62 ;
    RECT 57.145 75.86 58.06 76.62 ;
    RECT 58.54 75.86 59.46 76.62 ;
    RECT 59.94 75.86 60.16 76.62 ;
    RECT 60.64 75.86 60.855 76.62 ;
    RECT 61.335 75.86 61.555 76.62 ;
    RECT 62.035 75.86 62.25 76.62 ;
    RECT 62.73 75.86 63.65 76.62 ;
    RECT 64.13 75.86 64.345 76.62 ;
    RECT 64.825 75.86 65.045 76.62 ;
    RECT 65.525 75.86 65.745 76.62 ;
    RECT 66.225 75.86 66.445 76.62 ;
    RECT 66.925 75.86 67.14 76.62 ;
    RECT 67.62 75.86 67.84 76.62 ;
    RECT 68.32 75.86 69.235 76.62 ;
    RECT 69.715 75.86 69.935 76.62 ;
    RECT 70.415 75.86 70.635 76.62 ;
    RECT 71.115 75.86 71.335 76.62 ;
    RECT 71.815 75.86 72.035 76.62 ;
    RECT 72.515 75.86 72.735 76.62 ;
    RECT 73.215 75.86 73.435 76.62 ;
    RECT 73.915 75.86 74.835 76.62 ;
    RECT 75.315 75.86 75.535 76.62 ;
    RECT 76.015 75.86 76.225 76.62 ;
    RECT 76.705 75.86 76.92 76.62 ;
    RECT 77.4 75.86 77.62 76.62 ;
    RECT 78.1 75.86 78.32 76.62 ;
    RECT 78.8 75.86 79.02 76.62 ;
    RECT 79.5 75.86 81.115 76.62 ;
    RECT 81.595 75.86 81.815 76.62 ;
    RECT 82.295 75.86 82.515 76.62 ;
    RECT 82.995 75.86 83.055 76.62 ;
    RECT 83.055 75.77 83.335 76.71 ;
    RECT 83.335 75.86 83.505 76.62 ;
    RECT 26.71 75.1 26.88 75.86 ;
    RECT 26.88 75.01 27.16 75.95 ;
    RECT 27.16 75.1 27.32 75.86 ;
    RECT 27.8 75.1 28.02 75.86 ;
    RECT 28.5 75.1 28.72 75.86 ;
    RECT 29.2 75.1 30.815 75.86 ;
    RECT 31.295 75.1 31.515 75.86 ;
    RECT 31.995 75.1 32.21 75.86 ;
    RECT 32.69 75.1 32.91 75.86 ;
    RECT 33.39 75.1 33.61 75.86 ;
    RECT 34.09 75.1 34.31 75.86 ;
    RECT 34.79 75.1 35.005 75.86 ;
    RECT 35.485 75.1 36.405 75.86 ;
    RECT 36.885 75.1 37.105 75.86 ;
    RECT 37.585 75.1 37.8 75.86 ;
    RECT 38.28 75.1 38.5 75.86 ;
    RECT 38.98 75.1 39.2 75.86 ;
    RECT 39.68 75.1 39.895 75.86 ;
    RECT 40.375 75.1 40.595 75.86 ;
    RECT 41.075 75.1 41.995 75.86 ;
    RECT 42.475 75.1 42.69 75.86 ;
    RECT 43.17 75.1 43.39 75.86 ;
    RECT 43.87 75.1 44.09 75.86 ;
    RECT 44.57 75.1 44.79 75.86 ;
    RECT 45.27 75.1 45.485 75.86 ;
    RECT 45.965 75.1 46.185 75.86 ;
    RECT 46.665 75.1 47.58 75.86 ;
    RECT 48.06 75.1 48.28 75.86 ;
    RECT 48.76 75.1 48.98 75.86 ;
    RECT 49.46 75.1 49.68 75.86 ;
    RECT 50.16 75.1 50.375 75.86 ;
    RECT 50.855 75.1 51.775 75.86 ;
    RECT 52.255 75.1 53.17 75.86 ;
    RECT 53.65 75.1 53.87 75.86 ;
    RECT 54.35 75.1 54.57 75.86 ;
    RECT 55.05 75.1 55.265 75.86 ;
    RECT 55.745 75.1 55.965 75.86 ;
    RECT 56.445 75.1 56.665 75.86 ;
    RECT 57.145 75.1 58.06 75.86 ;
    RECT 58.54 75.1 59.46 75.86 ;
    RECT 59.94 75.1 60.16 75.86 ;
    RECT 60.64 75.1 60.855 75.86 ;
    RECT 61.335 75.1 61.555 75.86 ;
    RECT 62.035 75.1 62.25 75.86 ;
    RECT 62.73 75.1 63.65 75.86 ;
    RECT 64.13 75.1 64.345 75.86 ;
    RECT 64.825 75.1 65.045 75.86 ;
    RECT 65.525 75.1 65.745 75.86 ;
    RECT 66.225 75.1 66.445 75.86 ;
    RECT 66.925 75.1 67.14 75.86 ;
    RECT 67.62 75.1 67.84 75.86 ;
    RECT 68.32 75.1 69.235 75.86 ;
    RECT 69.715 75.1 69.935 75.86 ;
    RECT 70.415 75.1 70.635 75.86 ;
    RECT 71.115 75.1 71.335 75.86 ;
    RECT 71.815 75.1 72.035 75.86 ;
    RECT 72.515 75.1 72.735 75.86 ;
    RECT 73.215 75.1 73.435 75.86 ;
    RECT 73.915 75.1 74.835 75.86 ;
    RECT 75.315 75.1 75.535 75.86 ;
    RECT 76.015 75.1 76.225 75.86 ;
    RECT 76.705 75.1 76.92 75.86 ;
    RECT 77.4 75.1 77.62 75.86 ;
    RECT 78.1 75.1 78.32 75.86 ;
    RECT 78.8 75.1 79.02 75.86 ;
    RECT 79.5 75.1 81.115 75.86 ;
    RECT 81.595 75.1 81.815 75.86 ;
    RECT 82.295 75.1 82.515 75.86 ;
    RECT 82.995 75.1 83.055 75.86 ;
    RECT 83.055 75.01 83.335 75.95 ;
    RECT 83.335 75.1 83.505 75.86 ;
    RECT 26.71 74.34 26.88 75.1 ;
    RECT 26.88 74.25 27.16 75.19 ;
    RECT 27.16 74.34 27.32 75.1 ;
    RECT 27.8 74.34 28.02 75.1 ;
    RECT 28.5 74.34 28.72 75.1 ;
    RECT 29.2 74.34 30.815 75.1 ;
    RECT 31.295 74.34 31.515 75.1 ;
    RECT 31.995 74.34 32.21 75.1 ;
    RECT 32.69 74.34 32.91 75.1 ;
    RECT 33.39 74.34 33.61 75.1 ;
    RECT 34.09 74.34 34.31 75.1 ;
    RECT 34.79 74.34 35.005 75.1 ;
    RECT 35.485 74.34 36.405 75.1 ;
    RECT 36.885 74.34 37.105 75.1 ;
    RECT 37.585 74.34 37.8 75.1 ;
    RECT 38.28 74.34 38.5 75.1 ;
    RECT 38.98 74.34 39.2 75.1 ;
    RECT 39.68 74.34 39.895 75.1 ;
    RECT 40.375 74.34 40.595 75.1 ;
    RECT 41.075 74.34 41.995 75.1 ;
    RECT 42.475 74.34 42.69 75.1 ;
    RECT 43.17 74.34 43.39 75.1 ;
    RECT 43.87 74.34 44.09 75.1 ;
    RECT 44.57 74.34 44.79 75.1 ;
    RECT 45.27 74.34 45.485 75.1 ;
    RECT 45.965 74.34 46.185 75.1 ;
    RECT 46.665 74.34 47.58 75.1 ;
    RECT 48.06 74.34 48.28 75.1 ;
    RECT 48.76 74.34 48.98 75.1 ;
    RECT 49.46 74.34 49.68 75.1 ;
    RECT 50.16 74.34 50.375 75.1 ;
    RECT 50.855 74.34 51.775 75.1 ;
    RECT 52.255 74.34 53.17 75.1 ;
    RECT 53.65 74.34 53.87 75.1 ;
    RECT 54.35 74.34 54.57 75.1 ;
    RECT 55.05 74.34 55.265 75.1 ;
    RECT 55.745 74.34 55.965 75.1 ;
    RECT 56.445 74.34 56.665 75.1 ;
    RECT 57.145 74.34 58.06 75.1 ;
    RECT 58.54 74.34 59.46 75.1 ;
    RECT 59.94 74.34 60.16 75.1 ;
    RECT 60.64 74.34 60.855 75.1 ;
    RECT 61.335 74.34 61.555 75.1 ;
    RECT 62.035 74.34 62.25 75.1 ;
    RECT 62.73 74.34 63.65 75.1 ;
    RECT 64.13 74.34 64.345 75.1 ;
    RECT 64.825 74.34 65.045 75.1 ;
    RECT 65.525 74.34 65.745 75.1 ;
    RECT 66.225 74.34 66.445 75.1 ;
    RECT 66.925 74.34 67.14 75.1 ;
    RECT 67.62 74.34 67.84 75.1 ;
    RECT 68.32 74.34 69.235 75.1 ;
    RECT 69.715 74.34 69.935 75.1 ;
    RECT 70.415 74.34 70.635 75.1 ;
    RECT 71.115 74.34 71.335 75.1 ;
    RECT 71.815 74.34 72.035 75.1 ;
    RECT 72.515 74.34 72.735 75.1 ;
    RECT 73.215 74.34 73.435 75.1 ;
    RECT 73.915 74.34 74.835 75.1 ;
    RECT 75.315 74.34 75.535 75.1 ;
    RECT 76.015 74.34 76.225 75.1 ;
    RECT 76.705 74.34 76.92 75.1 ;
    RECT 77.4 74.34 77.62 75.1 ;
    RECT 78.1 74.34 78.32 75.1 ;
    RECT 78.8 74.34 79.02 75.1 ;
    RECT 79.5 74.34 81.115 75.1 ;
    RECT 81.595 74.34 81.815 75.1 ;
    RECT 82.295 74.34 82.515 75.1 ;
    RECT 82.995 74.34 83.055 75.1 ;
    RECT 83.055 74.25 83.335 75.19 ;
    RECT 83.335 74.34 83.505 75.1 ;
    RECT 26.71 73.58 26.88 74.34 ;
    RECT 26.88 73.49 27.16 74.43 ;
    RECT 27.16 73.58 27.32 74.34 ;
    RECT 27.8 73.58 28.02 74.34 ;
    RECT 28.5 73.58 28.72 74.34 ;
    RECT 29.2 73.58 30.815 74.34 ;
    RECT 31.295 73.58 31.515 74.34 ;
    RECT 31.995 73.58 32.21 74.34 ;
    RECT 32.69 73.58 32.91 74.34 ;
    RECT 33.39 73.58 33.61 74.34 ;
    RECT 34.09 73.58 34.31 74.34 ;
    RECT 34.79 73.58 35.005 74.34 ;
    RECT 35.485 73.58 36.405 74.34 ;
    RECT 36.885 73.58 37.105 74.34 ;
    RECT 37.585 73.58 37.8 74.34 ;
    RECT 38.28 73.58 38.5 74.34 ;
    RECT 38.98 73.58 39.2 74.34 ;
    RECT 39.68 73.58 39.895 74.34 ;
    RECT 40.375 73.58 40.595 74.34 ;
    RECT 41.075 73.58 41.995 74.34 ;
    RECT 42.475 73.58 42.69 74.34 ;
    RECT 43.17 73.58 43.39 74.34 ;
    RECT 43.87 73.58 44.09 74.34 ;
    RECT 44.57 73.58 44.79 74.34 ;
    RECT 45.27 73.58 45.485 74.34 ;
    RECT 45.965 73.58 46.185 74.34 ;
    RECT 46.665 73.58 47.58 74.34 ;
    RECT 48.06 73.58 48.28 74.34 ;
    RECT 48.76 73.58 48.98 74.34 ;
    RECT 49.46 73.58 49.68 74.34 ;
    RECT 50.16 73.58 50.375 74.34 ;
    RECT 50.855 73.58 51.775 74.34 ;
    RECT 52.255 73.58 53.17 74.34 ;
    RECT 53.65 73.58 53.87 74.34 ;
    RECT 54.35 73.58 54.57 74.34 ;
    RECT 55.05 73.58 55.265 74.34 ;
    RECT 55.745 73.58 55.965 74.34 ;
    RECT 56.445 73.58 56.665 74.34 ;
    RECT 57.145 73.58 58.06 74.34 ;
    RECT 58.54 73.58 59.46 74.34 ;
    RECT 59.94 73.58 60.16 74.34 ;
    RECT 60.64 73.58 60.855 74.34 ;
    RECT 61.335 73.58 61.555 74.34 ;
    RECT 62.035 73.58 62.25 74.34 ;
    RECT 62.73 73.58 63.65 74.34 ;
    RECT 64.13 73.58 64.345 74.34 ;
    RECT 64.825 73.58 65.045 74.34 ;
    RECT 65.525 73.58 65.745 74.34 ;
    RECT 66.225 73.58 66.445 74.34 ;
    RECT 66.925 73.58 67.14 74.34 ;
    RECT 67.62 73.58 67.84 74.34 ;
    RECT 68.32 73.58 69.235 74.34 ;
    RECT 69.715 73.58 69.935 74.34 ;
    RECT 70.415 73.58 70.635 74.34 ;
    RECT 71.115 73.58 71.335 74.34 ;
    RECT 71.815 73.58 72.035 74.34 ;
    RECT 72.515 73.58 72.735 74.34 ;
    RECT 73.215 73.58 73.435 74.34 ;
    RECT 73.915 73.58 74.835 74.34 ;
    RECT 75.315 73.58 75.535 74.34 ;
    RECT 76.015 73.58 76.225 74.34 ;
    RECT 76.705 73.58 76.92 74.34 ;
    RECT 77.4 73.58 77.62 74.34 ;
    RECT 78.1 73.58 78.32 74.34 ;
    RECT 78.8 73.58 79.02 74.34 ;
    RECT 79.5 73.58 81.115 74.34 ;
    RECT 81.595 73.58 81.815 74.34 ;
    RECT 82.295 73.58 82.515 74.34 ;
    RECT 82.995 73.58 83.055 74.34 ;
    RECT 83.055 73.49 83.335 74.43 ;
    RECT 83.335 73.58 83.505 74.34 ;
    RECT 26.71 72.82 26.88 73.58 ;
    RECT 26.88 72.73 27.16 73.67 ;
    RECT 27.16 72.82 27.32 73.58 ;
    RECT 27.8 72.82 28.02 73.58 ;
    RECT 28.5 72.82 28.72 73.58 ;
    RECT 29.2 72.82 30.815 73.58 ;
    RECT 31.295 72.82 31.515 73.58 ;
    RECT 31.995 72.82 32.21 73.58 ;
    RECT 32.69 72.82 32.91 73.58 ;
    RECT 33.39 72.82 33.61 73.58 ;
    RECT 34.09 72.82 34.31 73.58 ;
    RECT 34.79 72.82 35.005 73.58 ;
    RECT 35.485 72.82 36.405 73.58 ;
    RECT 36.885 72.82 37.105 73.58 ;
    RECT 37.585 72.82 37.8 73.58 ;
    RECT 38.28 72.82 38.5 73.58 ;
    RECT 38.98 72.82 39.2 73.58 ;
    RECT 39.68 72.82 39.895 73.58 ;
    RECT 40.375 72.82 40.595 73.58 ;
    RECT 41.075 72.82 41.995 73.58 ;
    RECT 42.475 72.82 42.69 73.58 ;
    RECT 43.17 72.82 43.39 73.58 ;
    RECT 43.87 72.82 44.09 73.58 ;
    RECT 44.57 72.82 44.79 73.58 ;
    RECT 45.27 72.82 45.485 73.58 ;
    RECT 45.965 72.82 46.185 73.58 ;
    RECT 46.665 72.82 47.58 73.58 ;
    RECT 48.06 72.82 48.28 73.58 ;
    RECT 48.76 72.82 48.98 73.58 ;
    RECT 49.46 72.82 49.68 73.58 ;
    RECT 50.16 72.82 50.375 73.58 ;
    RECT 50.855 72.82 51.775 73.58 ;
    RECT 52.255 72.82 53.17 73.58 ;
    RECT 53.65 72.82 53.87 73.58 ;
    RECT 54.35 72.82 54.57 73.58 ;
    RECT 55.05 72.82 55.265 73.58 ;
    RECT 55.745 72.82 55.965 73.58 ;
    RECT 56.445 72.82 56.665 73.58 ;
    RECT 57.145 72.82 58.06 73.58 ;
    RECT 58.54 72.82 59.46 73.58 ;
    RECT 59.94 72.82 60.16 73.58 ;
    RECT 60.64 72.82 60.855 73.58 ;
    RECT 61.335 72.82 61.555 73.58 ;
    RECT 62.035 72.82 62.25 73.58 ;
    RECT 62.73 72.82 63.65 73.58 ;
    RECT 64.13 72.82 64.345 73.58 ;
    RECT 64.825 72.82 65.045 73.58 ;
    RECT 65.525 72.82 65.745 73.58 ;
    RECT 66.225 72.82 66.445 73.58 ;
    RECT 66.925 72.82 67.14 73.58 ;
    RECT 67.62 72.82 67.84 73.58 ;
    RECT 68.32 72.82 69.235 73.58 ;
    RECT 69.715 72.82 69.935 73.58 ;
    RECT 70.415 72.82 70.635 73.58 ;
    RECT 71.115 72.82 71.335 73.58 ;
    RECT 71.815 72.82 72.035 73.58 ;
    RECT 72.515 72.82 72.735 73.58 ;
    RECT 73.215 72.82 73.435 73.58 ;
    RECT 73.915 72.82 74.835 73.58 ;
    RECT 75.315 72.82 75.535 73.58 ;
    RECT 76.015 72.82 76.225 73.58 ;
    RECT 76.705 72.82 76.92 73.58 ;
    RECT 77.4 72.82 77.62 73.58 ;
    RECT 78.1 72.82 78.32 73.58 ;
    RECT 78.8 72.82 79.02 73.58 ;
    RECT 79.5 72.82 81.115 73.58 ;
    RECT 81.595 72.82 81.815 73.58 ;
    RECT 82.295 72.82 82.515 73.58 ;
    RECT 82.995 72.82 83.055 73.58 ;
    RECT 83.055 72.73 83.335 73.67 ;
    RECT 83.335 72.82 83.505 73.58 ;
    RECT 26.71 72.06 26.88 72.82 ;
    RECT 26.88 71.97 27.16 72.91 ;
    RECT 27.16 72.06 27.32 72.82 ;
    RECT 27.8 72.06 28.02 72.82 ;
    RECT 28.5 72.06 28.72 72.82 ;
    RECT 29.2 72.06 30.815 72.82 ;
    RECT 31.295 72.06 31.515 72.82 ;
    RECT 31.995 72.06 32.21 72.82 ;
    RECT 32.69 72.06 32.91 72.82 ;
    RECT 33.39 72.06 33.61 72.82 ;
    RECT 34.09 72.06 34.31 72.82 ;
    RECT 34.79 72.06 35.005 72.82 ;
    RECT 35.485 72.06 36.405 72.82 ;
    RECT 36.885 72.06 37.105 72.82 ;
    RECT 37.585 72.06 37.8 72.82 ;
    RECT 38.28 72.06 38.5 72.82 ;
    RECT 38.98 72.06 39.2 72.82 ;
    RECT 39.68 72.06 39.895 72.82 ;
    RECT 40.375 72.06 40.595 72.82 ;
    RECT 41.075 72.06 41.995 72.82 ;
    RECT 42.475 72.06 42.69 72.82 ;
    RECT 43.17 72.06 43.39 72.82 ;
    RECT 43.87 72.06 44.09 72.82 ;
    RECT 44.57 72.06 44.79 72.82 ;
    RECT 45.27 72.06 45.485 72.82 ;
    RECT 45.965 72.06 46.185 72.82 ;
    RECT 46.665 72.06 47.58 72.82 ;
    RECT 48.06 72.06 48.28 72.82 ;
    RECT 48.76 72.06 48.98 72.82 ;
    RECT 49.46 72.06 49.68 72.82 ;
    RECT 50.16 72.06 50.375 72.82 ;
    RECT 50.855 72.06 51.775 72.82 ;
    RECT 52.255 72.06 53.17 72.82 ;
    RECT 53.65 72.06 53.87 72.82 ;
    RECT 54.35 72.06 54.57 72.82 ;
    RECT 55.05 72.06 55.265 72.82 ;
    RECT 55.745 72.06 55.965 72.82 ;
    RECT 56.445 72.06 56.665 72.82 ;
    RECT 57.145 72.06 58.06 72.82 ;
    RECT 58.54 72.06 59.46 72.82 ;
    RECT 59.94 72.06 60.16 72.82 ;
    RECT 60.64 72.06 60.855 72.82 ;
    RECT 61.335 72.06 61.555 72.82 ;
    RECT 62.035 72.06 62.25 72.82 ;
    RECT 62.73 72.06 63.65 72.82 ;
    RECT 64.13 72.06 64.345 72.82 ;
    RECT 64.825 72.06 65.045 72.82 ;
    RECT 65.525 72.06 65.745 72.82 ;
    RECT 66.225 72.06 66.445 72.82 ;
    RECT 66.925 72.06 67.14 72.82 ;
    RECT 67.62 72.06 67.84 72.82 ;
    RECT 68.32 72.06 69.235 72.82 ;
    RECT 69.715 72.06 69.935 72.82 ;
    RECT 70.415 72.06 70.635 72.82 ;
    RECT 71.115 72.06 71.335 72.82 ;
    RECT 71.815 72.06 72.035 72.82 ;
    RECT 72.515 72.06 72.735 72.82 ;
    RECT 73.215 72.06 73.435 72.82 ;
    RECT 73.915 72.06 74.835 72.82 ;
    RECT 75.315 72.06 75.535 72.82 ;
    RECT 76.015 72.06 76.225 72.82 ;
    RECT 76.705 72.06 76.92 72.82 ;
    RECT 77.4 72.06 77.62 72.82 ;
    RECT 78.1 72.06 78.32 72.82 ;
    RECT 78.8 72.06 79.02 72.82 ;
    RECT 79.5 72.06 81.115 72.82 ;
    RECT 81.595 72.06 81.815 72.82 ;
    RECT 82.295 72.06 82.515 72.82 ;
    RECT 82.995 72.06 83.055 72.82 ;
    RECT 83.055 71.97 83.335 72.91 ;
    RECT 83.335 72.06 83.505 72.82 ;
    RECT 26.71 71.3 26.88 72.06 ;
    RECT 26.88 71.21 27.16 72.15 ;
    RECT 27.16 71.3 27.32 72.06 ;
    RECT 27.8 71.3 28.02 72.06 ;
    RECT 28.5 71.3 28.72 72.06 ;
    RECT 29.2 71.3 30.815 72.06 ;
    RECT 31.295 71.3 31.515 72.06 ;
    RECT 31.995 71.3 32.21 72.06 ;
    RECT 32.69 71.3 32.91 72.06 ;
    RECT 33.39 71.3 33.61 72.06 ;
    RECT 34.09 71.3 34.31 72.06 ;
    RECT 34.79 71.3 35.005 72.06 ;
    RECT 35.485 71.3 36.405 72.06 ;
    RECT 36.885 71.3 37.105 72.06 ;
    RECT 37.585 71.3 37.8 72.06 ;
    RECT 38.28 71.3 38.5 72.06 ;
    RECT 38.98 71.3 39.2 72.06 ;
    RECT 39.68 71.3 39.895 72.06 ;
    RECT 40.375 71.3 40.595 72.06 ;
    RECT 41.075 71.3 41.995 72.06 ;
    RECT 42.475 71.3 42.69 72.06 ;
    RECT 43.17 71.3 43.39 72.06 ;
    RECT 43.87 71.3 44.09 72.06 ;
    RECT 44.57 71.3 44.79 72.06 ;
    RECT 45.27 71.3 45.485 72.06 ;
    RECT 45.965 71.3 46.185 72.06 ;
    RECT 46.665 71.3 47.58 72.06 ;
    RECT 48.06 71.3 48.28 72.06 ;
    RECT 48.76 71.3 48.98 72.06 ;
    RECT 49.46 71.3 49.68 72.06 ;
    RECT 50.16 71.3 50.375 72.06 ;
    RECT 50.855 71.3 51.775 72.06 ;
    RECT 52.255 71.3 53.17 72.06 ;
    RECT 53.65 71.3 53.87 72.06 ;
    RECT 54.35 71.3 54.57 72.06 ;
    RECT 55.05 71.3 55.265 72.06 ;
    RECT 55.745 71.3 55.965 72.06 ;
    RECT 56.445 71.3 56.665 72.06 ;
    RECT 57.145 71.3 58.06 72.06 ;
    RECT 58.54 71.3 59.46 72.06 ;
    RECT 59.94 71.3 60.16 72.06 ;
    RECT 60.64 71.3 60.855 72.06 ;
    RECT 61.335 71.3 61.555 72.06 ;
    RECT 62.035 71.3 62.25 72.06 ;
    RECT 62.73 71.3 63.65 72.06 ;
    RECT 64.13 71.3 64.345 72.06 ;
    RECT 64.825 71.3 65.045 72.06 ;
    RECT 65.525 71.3 65.745 72.06 ;
    RECT 66.225 71.3 66.445 72.06 ;
    RECT 66.925 71.3 67.14 72.06 ;
    RECT 67.62 71.3 67.84 72.06 ;
    RECT 68.32 71.3 69.235 72.06 ;
    RECT 69.715 71.3 69.935 72.06 ;
    RECT 70.415 71.3 70.635 72.06 ;
    RECT 71.115 71.3 71.335 72.06 ;
    RECT 71.815 71.3 72.035 72.06 ;
    RECT 72.515 71.3 72.735 72.06 ;
    RECT 73.215 71.3 73.435 72.06 ;
    RECT 73.915 71.3 74.835 72.06 ;
    RECT 75.315 71.3 75.535 72.06 ;
    RECT 76.015 71.3 76.225 72.06 ;
    RECT 76.705 71.3 76.92 72.06 ;
    RECT 77.4 71.3 77.62 72.06 ;
    RECT 78.1 71.3 78.32 72.06 ;
    RECT 78.8 71.3 79.02 72.06 ;
    RECT 79.5 71.3 81.115 72.06 ;
    RECT 81.595 71.3 81.815 72.06 ;
    RECT 82.295 71.3 82.515 72.06 ;
    RECT 82.995 71.3 83.055 72.06 ;
    RECT 83.055 71.21 83.335 72.15 ;
    RECT 83.335 71.3 83.505 72.06 ;
    RECT 26.71 70.54 26.88 71.3 ;
    RECT 26.88 70.45 27.16 71.39 ;
    RECT 27.16 70.54 27.32 71.3 ;
    RECT 27.8 70.54 28.02 71.3 ;
    RECT 28.5 70.54 28.72 71.3 ;
    RECT 29.2 70.54 30.815 71.3 ;
    RECT 31.295 70.54 31.515 71.3 ;
    RECT 31.995 70.54 32.21 71.3 ;
    RECT 32.69 70.54 32.91 71.3 ;
    RECT 33.39 70.54 33.61 71.3 ;
    RECT 34.09 70.54 34.31 71.3 ;
    RECT 34.79 70.54 35.005 71.3 ;
    RECT 35.485 70.54 36.405 71.3 ;
    RECT 36.885 70.54 37.105 71.3 ;
    RECT 37.585 70.54 37.8 71.3 ;
    RECT 38.28 70.54 38.5 71.3 ;
    RECT 38.98 70.54 39.2 71.3 ;
    RECT 39.68 70.54 39.895 71.3 ;
    RECT 40.375 70.54 40.595 71.3 ;
    RECT 41.075 70.54 41.995 71.3 ;
    RECT 42.475 70.54 42.69 71.3 ;
    RECT 43.17 70.54 43.39 71.3 ;
    RECT 43.87 70.54 44.09 71.3 ;
    RECT 44.57 70.54 44.79 71.3 ;
    RECT 45.27 70.54 45.485 71.3 ;
    RECT 45.965 70.54 46.185 71.3 ;
    RECT 46.665 70.54 47.58 71.3 ;
    RECT 48.06 70.54 48.28 71.3 ;
    RECT 48.76 70.54 48.98 71.3 ;
    RECT 49.46 70.54 49.68 71.3 ;
    RECT 50.16 70.54 50.375 71.3 ;
    RECT 50.855 70.54 51.775 71.3 ;
    RECT 52.255 70.54 53.17 71.3 ;
    RECT 53.65 70.54 53.87 71.3 ;
    RECT 54.35 70.54 54.57 71.3 ;
    RECT 55.05 70.54 55.265 71.3 ;
    RECT 55.745 70.54 55.965 71.3 ;
    RECT 56.445 70.54 56.665 71.3 ;
    RECT 57.145 70.54 58.06 71.3 ;
    RECT 58.54 70.54 59.46 71.3 ;
    RECT 59.94 70.54 60.16 71.3 ;
    RECT 60.64 70.54 60.855 71.3 ;
    RECT 61.335 70.54 61.555 71.3 ;
    RECT 62.035 70.54 62.25 71.3 ;
    RECT 62.73 70.54 63.65 71.3 ;
    RECT 64.13 70.54 64.345 71.3 ;
    RECT 64.825 70.54 65.045 71.3 ;
    RECT 65.525 70.54 65.745 71.3 ;
    RECT 66.225 70.54 66.445 71.3 ;
    RECT 66.925 70.54 67.14 71.3 ;
    RECT 67.62 70.54 67.84 71.3 ;
    RECT 68.32 70.54 69.235 71.3 ;
    RECT 69.715 70.54 69.935 71.3 ;
    RECT 70.415 70.54 70.635 71.3 ;
    RECT 71.115 70.54 71.335 71.3 ;
    RECT 71.815 70.54 72.035 71.3 ;
    RECT 72.515 70.54 72.735 71.3 ;
    RECT 73.215 70.54 73.435 71.3 ;
    RECT 73.915 70.54 74.835 71.3 ;
    RECT 75.315 70.54 75.535 71.3 ;
    RECT 76.015 70.54 76.225 71.3 ;
    RECT 76.705 70.54 76.92 71.3 ;
    RECT 77.4 70.54 77.62 71.3 ;
    RECT 78.1 70.54 78.32 71.3 ;
    RECT 78.8 70.54 79.02 71.3 ;
    RECT 79.5 70.54 81.115 71.3 ;
    RECT 81.595 70.54 81.815 71.3 ;
    RECT 82.295 70.54 82.515 71.3 ;
    RECT 82.995 70.54 83.055 71.3 ;
    RECT 83.055 70.45 83.335 71.39 ;
    RECT 83.335 70.54 83.505 71.3 ;
    RECT 26.71 69.78 26.88 70.54 ;
    RECT 26.88 69.69 27.16 70.63 ;
    RECT 27.16 69.78 27.32 70.54 ;
    RECT 27.8 69.78 28.02 70.54 ;
    RECT 28.5 69.78 28.72 70.54 ;
    RECT 29.2 69.78 30.815 70.54 ;
    RECT 31.295 69.78 31.515 70.54 ;
    RECT 31.995 69.78 32.21 70.54 ;
    RECT 32.69 69.78 32.91 70.54 ;
    RECT 33.39 69.78 33.61 70.54 ;
    RECT 34.09 69.78 34.31 70.54 ;
    RECT 34.79 69.78 35.005 70.54 ;
    RECT 35.485 69.78 36.405 70.54 ;
    RECT 36.885 69.78 37.105 70.54 ;
    RECT 37.585 69.78 37.8 70.54 ;
    RECT 38.28 69.78 38.5 70.54 ;
    RECT 38.98 69.78 39.2 70.54 ;
    RECT 39.68 69.78 39.895 70.54 ;
    RECT 40.375 69.78 40.595 70.54 ;
    RECT 41.075 69.78 41.995 70.54 ;
    RECT 42.475 69.78 42.69 70.54 ;
    RECT 43.17 69.78 43.39 70.54 ;
    RECT 43.87 69.78 44.09 70.54 ;
    RECT 44.57 69.78 44.79 70.54 ;
    RECT 45.27 69.78 45.485 70.54 ;
    RECT 45.965 69.78 46.185 70.54 ;
    RECT 46.665 69.78 47.58 70.54 ;
    RECT 48.06 69.78 48.28 70.54 ;
    RECT 48.76 69.78 48.98 70.54 ;
    RECT 49.46 69.78 49.68 70.54 ;
    RECT 50.16 69.78 50.375 70.54 ;
    RECT 50.855 69.78 51.775 70.54 ;
    RECT 52.255 69.78 53.17 70.54 ;
    RECT 53.65 69.78 53.87 70.54 ;
    RECT 54.35 69.78 54.57 70.54 ;
    RECT 55.05 69.78 55.265 70.54 ;
    RECT 55.745 69.78 55.965 70.54 ;
    RECT 56.445 69.78 56.665 70.54 ;
    RECT 57.145 69.78 58.06 70.54 ;
    RECT 58.54 69.78 59.46 70.54 ;
    RECT 59.94 69.78 60.16 70.54 ;
    RECT 60.64 69.78 60.855 70.54 ;
    RECT 61.335 69.78 61.555 70.54 ;
    RECT 62.035 69.78 62.25 70.54 ;
    RECT 62.73 69.78 63.65 70.54 ;
    RECT 64.13 69.78 64.345 70.54 ;
    RECT 64.825 69.78 65.045 70.54 ;
    RECT 65.525 69.78 65.745 70.54 ;
    RECT 66.225 69.78 66.445 70.54 ;
    RECT 66.925 69.78 67.14 70.54 ;
    RECT 67.62 69.78 67.84 70.54 ;
    RECT 68.32 69.78 69.235 70.54 ;
    RECT 69.715 69.78 69.935 70.54 ;
    RECT 70.415 69.78 70.635 70.54 ;
    RECT 71.115 69.78 71.335 70.54 ;
    RECT 71.815 69.78 72.035 70.54 ;
    RECT 72.515 69.78 72.735 70.54 ;
    RECT 73.215 69.78 73.435 70.54 ;
    RECT 73.915 69.78 74.835 70.54 ;
    RECT 75.315 69.78 75.535 70.54 ;
    RECT 76.015 69.78 76.225 70.54 ;
    RECT 76.705 69.78 76.92 70.54 ;
    RECT 77.4 69.78 77.62 70.54 ;
    RECT 78.1 69.78 78.32 70.54 ;
    RECT 78.8 69.78 79.02 70.54 ;
    RECT 79.5 69.78 81.115 70.54 ;
    RECT 81.595 69.78 81.815 70.54 ;
    RECT 82.295 69.78 82.515 70.54 ;
    RECT 82.995 69.78 83.055 70.54 ;
    RECT 83.055 69.69 83.335 70.63 ;
    RECT 83.335 69.78 83.505 70.54 ;
    RECT 26.71 69.02 26.88 69.78 ;
    RECT 26.88 68.93 27.16 69.87 ;
    RECT 27.16 69.02 27.32 69.78 ;
    RECT 27.8 69.02 28.02 69.78 ;
    RECT 28.5 69.02 28.72 69.78 ;
    RECT 29.2 69.02 30.815 69.78 ;
    RECT 31.295 69.02 31.515 69.78 ;
    RECT 31.995 69.02 32.21 69.78 ;
    RECT 32.69 69.02 32.91 69.78 ;
    RECT 33.39 69.02 33.61 69.78 ;
    RECT 34.09 69.02 34.31 69.78 ;
    RECT 34.79 69.02 35.005 69.78 ;
    RECT 35.485 69.02 36.405 69.78 ;
    RECT 36.885 69.02 37.105 69.78 ;
    RECT 37.585 69.02 37.8 69.78 ;
    RECT 38.28 69.02 38.5 69.78 ;
    RECT 38.98 69.02 39.2 69.78 ;
    RECT 39.68 69.02 39.895 69.78 ;
    RECT 40.375 69.02 40.595 69.78 ;
    RECT 41.075 69.02 41.995 69.78 ;
    RECT 42.475 69.02 42.69 69.78 ;
    RECT 43.17 69.02 43.39 69.78 ;
    RECT 43.87 69.02 44.09 69.78 ;
    RECT 44.57 69.02 44.79 69.78 ;
    RECT 45.27 69.02 45.485 69.78 ;
    RECT 45.965 69.02 46.185 69.78 ;
    RECT 46.665 69.02 47.58 69.78 ;
    RECT 48.06 69.02 48.28 69.78 ;
    RECT 48.76 69.02 48.98 69.78 ;
    RECT 49.46 69.02 49.68 69.78 ;
    RECT 50.16 69.02 50.375 69.78 ;
    RECT 50.855 69.02 51.775 69.78 ;
    RECT 52.255 69.02 53.17 69.78 ;
    RECT 53.65 69.02 53.87 69.78 ;
    RECT 54.35 69.02 54.57 69.78 ;
    RECT 55.05 69.02 55.265 69.78 ;
    RECT 55.745 69.02 55.965 69.78 ;
    RECT 56.445 69.02 56.665 69.78 ;
    RECT 57.145 69.02 58.06 69.78 ;
    RECT 58.54 69.02 59.46 69.78 ;
    RECT 59.94 69.02 60.16 69.78 ;
    RECT 60.64 69.02 60.855 69.78 ;
    RECT 61.335 69.02 61.555 69.78 ;
    RECT 62.035 69.02 62.25 69.78 ;
    RECT 62.73 69.02 63.65 69.78 ;
    RECT 64.13 69.02 64.345 69.78 ;
    RECT 64.825 69.02 65.045 69.78 ;
    RECT 65.525 69.02 65.745 69.78 ;
    RECT 66.225 69.02 66.445 69.78 ;
    RECT 66.925 69.02 67.14 69.78 ;
    RECT 67.62 69.02 67.84 69.78 ;
    RECT 68.32 69.02 69.235 69.78 ;
    RECT 69.715 69.02 69.935 69.78 ;
    RECT 70.415 69.02 70.635 69.78 ;
    RECT 71.115 69.02 71.335 69.78 ;
    RECT 71.815 69.02 72.035 69.78 ;
    RECT 72.515 69.02 72.735 69.78 ;
    RECT 73.215 69.02 73.435 69.78 ;
    RECT 73.915 69.02 74.835 69.78 ;
    RECT 75.315 69.02 75.535 69.78 ;
    RECT 76.015 69.02 76.225 69.78 ;
    RECT 76.705 69.02 76.92 69.78 ;
    RECT 77.4 69.02 77.62 69.78 ;
    RECT 78.1 69.02 78.32 69.78 ;
    RECT 78.8 69.02 79.02 69.78 ;
    RECT 79.5 69.02 81.115 69.78 ;
    RECT 81.595 69.02 81.815 69.78 ;
    RECT 82.295 69.02 82.515 69.78 ;
    RECT 82.995 69.02 83.055 69.78 ;
    RECT 83.055 68.93 83.335 69.87 ;
    RECT 83.335 69.02 83.505 69.78 ;
    RECT 26.71 68.26 26.88 69.02 ;
    RECT 26.88 68.17 27.16 69.11 ;
    RECT 27.16 68.26 27.32 69.02 ;
    RECT 27.8 68.26 28.02 69.02 ;
    RECT 28.5 68.26 28.72 69.02 ;
    RECT 29.2 68.26 30.815 69.02 ;
    RECT 31.295 68.26 31.515 69.02 ;
    RECT 31.995 68.26 32.21 69.02 ;
    RECT 32.69 68.26 32.91 69.02 ;
    RECT 33.39 68.26 33.61 69.02 ;
    RECT 34.09 68.26 34.31 69.02 ;
    RECT 34.79 68.26 35.005 69.02 ;
    RECT 35.485 68.26 36.405 69.02 ;
    RECT 36.885 68.26 37.105 69.02 ;
    RECT 37.585 68.26 37.8 69.02 ;
    RECT 38.28 68.26 38.5 69.02 ;
    RECT 38.98 68.26 39.2 69.02 ;
    RECT 39.68 68.26 39.895 69.02 ;
    RECT 40.375 68.26 40.595 69.02 ;
    RECT 41.075 68.26 41.995 69.02 ;
    RECT 42.475 68.26 42.69 69.02 ;
    RECT 43.17 68.26 43.39 69.02 ;
    RECT 43.87 68.26 44.09 69.02 ;
    RECT 44.57 68.26 44.79 69.02 ;
    RECT 45.27 68.26 45.485 69.02 ;
    RECT 45.965 68.26 46.185 69.02 ;
    RECT 46.665 68.26 47.58 69.02 ;
    RECT 48.06 68.26 48.28 69.02 ;
    RECT 48.76 68.26 48.98 69.02 ;
    RECT 49.46 68.26 49.68 69.02 ;
    RECT 50.16 68.26 50.375 69.02 ;
    RECT 50.855 68.26 51.775 69.02 ;
    RECT 52.255 68.26 53.17 69.02 ;
    RECT 53.65 68.26 53.87 69.02 ;
    RECT 54.35 68.26 54.57 69.02 ;
    RECT 55.05 68.26 55.265 69.02 ;
    RECT 55.745 68.26 55.965 69.02 ;
    RECT 56.445 68.26 56.665 69.02 ;
    RECT 57.145 68.26 58.06 69.02 ;
    RECT 58.54 68.26 59.46 69.02 ;
    RECT 59.94 68.26 60.16 69.02 ;
    RECT 60.64 68.26 60.855 69.02 ;
    RECT 61.335 68.26 61.555 69.02 ;
    RECT 62.035 68.26 62.25 69.02 ;
    RECT 62.73 68.26 63.65 69.02 ;
    RECT 64.13 68.26 64.345 69.02 ;
    RECT 64.825 68.26 65.045 69.02 ;
    RECT 65.525 68.26 65.745 69.02 ;
    RECT 66.225 68.26 66.445 69.02 ;
    RECT 66.925 68.26 67.14 69.02 ;
    RECT 67.62 68.26 67.84 69.02 ;
    RECT 68.32 68.26 69.235 69.02 ;
    RECT 69.715 68.26 69.935 69.02 ;
    RECT 70.415 68.26 70.635 69.02 ;
    RECT 71.115 68.26 71.335 69.02 ;
    RECT 71.815 68.26 72.035 69.02 ;
    RECT 72.515 68.26 72.735 69.02 ;
    RECT 73.215 68.26 73.435 69.02 ;
    RECT 73.915 68.26 74.835 69.02 ;
    RECT 75.315 68.26 75.535 69.02 ;
    RECT 76.015 68.26 76.225 69.02 ;
    RECT 76.705 68.26 76.92 69.02 ;
    RECT 77.4 68.26 77.62 69.02 ;
    RECT 78.1 68.26 78.32 69.02 ;
    RECT 78.8 68.26 79.02 69.02 ;
    RECT 79.5 68.26 81.115 69.02 ;
    RECT 81.595 68.26 81.815 69.02 ;
    RECT 82.295 68.26 82.515 69.02 ;
    RECT 82.995 68.26 83.055 69.02 ;
    RECT 83.055 68.17 83.335 69.11 ;
    RECT 83.335 68.26 83.505 69.02 ;
    RECT 26.71 67.5 26.88 68.26 ;
    RECT 26.88 67.41 27.16 68.35 ;
    RECT 27.16 67.5 27.32 68.26 ;
    RECT 27.8 67.5 28.02 68.26 ;
    RECT 28.5 67.5 28.72 68.26 ;
    RECT 29.2 67.5 30.815 68.26 ;
    RECT 31.295 67.5 31.515 68.26 ;
    RECT 31.995 67.5 32.21 68.26 ;
    RECT 32.69 67.5 32.91 68.26 ;
    RECT 33.39 67.5 33.61 68.26 ;
    RECT 34.09 67.5 34.31 68.26 ;
    RECT 34.79 67.5 35.005 68.26 ;
    RECT 35.485 67.5 36.405 68.26 ;
    RECT 36.885 67.5 37.105 68.26 ;
    RECT 37.585 67.5 37.8 68.26 ;
    RECT 38.28 67.5 38.5 68.26 ;
    RECT 38.98 67.5 39.2 68.26 ;
    RECT 39.68 67.5 39.895 68.26 ;
    RECT 40.375 67.5 40.595 68.26 ;
    RECT 41.075 67.5 41.995 68.26 ;
    RECT 42.475 67.5 42.69 68.26 ;
    RECT 43.17 67.5 43.39 68.26 ;
    RECT 43.87 67.5 44.09 68.26 ;
    RECT 44.57 67.5 44.79 68.26 ;
    RECT 45.27 67.5 45.485 68.26 ;
    RECT 45.965 67.5 46.185 68.26 ;
    RECT 46.665 67.5 47.58 68.26 ;
    RECT 48.06 67.5 48.28 68.26 ;
    RECT 48.76 67.5 48.98 68.26 ;
    RECT 49.46 67.5 49.68 68.26 ;
    RECT 50.16 67.5 50.375 68.26 ;
    RECT 50.855 67.5 51.775 68.26 ;
    RECT 52.255 67.5 53.17 68.26 ;
    RECT 53.65 67.5 53.87 68.26 ;
    RECT 54.35 67.5 54.57 68.26 ;
    RECT 55.05 67.5 55.265 68.26 ;
    RECT 55.745 67.5 55.965 68.26 ;
    RECT 56.445 67.5 56.665 68.26 ;
    RECT 57.145 67.5 58.06 68.26 ;
    RECT 58.54 67.5 59.46 68.26 ;
    RECT 59.94 67.5 60.16 68.26 ;
    RECT 60.64 67.5 60.855 68.26 ;
    RECT 61.335 67.5 61.555 68.26 ;
    RECT 62.035 67.5 62.25 68.26 ;
    RECT 62.73 67.5 63.65 68.26 ;
    RECT 64.13 67.5 64.345 68.26 ;
    RECT 64.825 67.5 65.045 68.26 ;
    RECT 65.525 67.5 65.745 68.26 ;
    RECT 66.225 67.5 66.445 68.26 ;
    RECT 66.925 67.5 67.14 68.26 ;
    RECT 67.62 67.5 67.84 68.26 ;
    RECT 68.32 67.5 69.235 68.26 ;
    RECT 69.715 67.5 69.935 68.26 ;
    RECT 70.415 67.5 70.635 68.26 ;
    RECT 71.115 67.5 71.335 68.26 ;
    RECT 71.815 67.5 72.035 68.26 ;
    RECT 72.515 67.5 72.735 68.26 ;
    RECT 73.215 67.5 73.435 68.26 ;
    RECT 73.915 67.5 74.835 68.26 ;
    RECT 75.315 67.5 75.535 68.26 ;
    RECT 76.015 67.5 76.225 68.26 ;
    RECT 76.705 67.5 76.92 68.26 ;
    RECT 77.4 67.5 77.62 68.26 ;
    RECT 78.1 67.5 78.32 68.26 ;
    RECT 78.8 67.5 79.02 68.26 ;
    RECT 79.5 67.5 81.115 68.26 ;
    RECT 81.595 67.5 81.815 68.26 ;
    RECT 82.295 67.5 82.515 68.26 ;
    RECT 82.995 67.5 83.055 68.26 ;
    RECT 83.055 67.41 83.335 68.35 ;
    RECT 83.335 67.5 83.505 68.26 ;
    RECT 26.71 66.74 26.88 67.5 ;
    RECT 26.88 66.65 27.16 67.59 ;
    RECT 27.16 66.74 27.32 67.5 ;
    RECT 27.8 66.74 28.02 67.5 ;
    RECT 28.5 66.74 28.72 67.5 ;
    RECT 29.2 66.74 30.815 67.5 ;
    RECT 31.295 66.74 31.515 67.5 ;
    RECT 31.995 66.74 32.21 67.5 ;
    RECT 32.69 66.74 32.91 67.5 ;
    RECT 33.39 66.74 33.61 67.5 ;
    RECT 34.09 66.74 34.31 67.5 ;
    RECT 34.79 66.74 35.005 67.5 ;
    RECT 35.485 66.74 36.405 67.5 ;
    RECT 36.885 66.74 37.105 67.5 ;
    RECT 37.585 66.74 37.8 67.5 ;
    RECT 38.28 66.74 38.5 67.5 ;
    RECT 38.98 66.74 39.2 67.5 ;
    RECT 39.68 66.74 39.895 67.5 ;
    RECT 40.375 66.74 40.595 67.5 ;
    RECT 41.075 66.74 41.995 67.5 ;
    RECT 42.475 66.74 42.69 67.5 ;
    RECT 43.17 66.74 43.39 67.5 ;
    RECT 43.87 66.74 44.09 67.5 ;
    RECT 44.57 66.74 44.79 67.5 ;
    RECT 45.27 66.74 45.485 67.5 ;
    RECT 45.965 66.74 46.185 67.5 ;
    RECT 46.665 66.74 47.58 67.5 ;
    RECT 48.06 66.74 48.28 67.5 ;
    RECT 48.76 66.74 48.98 67.5 ;
    RECT 49.46 66.74 49.68 67.5 ;
    RECT 50.16 66.74 50.375 67.5 ;
    RECT 50.855 66.74 51.775 67.5 ;
    RECT 52.255 66.74 53.17 67.5 ;
    RECT 53.65 66.74 53.87 67.5 ;
    RECT 54.35 66.74 54.57 67.5 ;
    RECT 55.05 66.74 55.265 67.5 ;
    RECT 55.745 66.74 55.965 67.5 ;
    RECT 56.445 66.74 56.665 67.5 ;
    RECT 57.145 66.74 58.06 67.5 ;
    RECT 58.54 66.74 59.46 67.5 ;
    RECT 59.94 66.74 60.16 67.5 ;
    RECT 60.64 66.74 60.855 67.5 ;
    RECT 61.335 66.74 61.555 67.5 ;
    RECT 62.035 66.74 62.25 67.5 ;
    RECT 62.73 66.74 63.65 67.5 ;
    RECT 64.13 66.74 64.345 67.5 ;
    RECT 64.825 66.74 65.045 67.5 ;
    RECT 65.525 66.74 65.745 67.5 ;
    RECT 66.225 66.74 66.445 67.5 ;
    RECT 66.925 66.74 67.14 67.5 ;
    RECT 67.62 66.74 67.84 67.5 ;
    RECT 68.32 66.74 69.235 67.5 ;
    RECT 69.715 66.74 69.935 67.5 ;
    RECT 70.415 66.74 70.635 67.5 ;
    RECT 71.115 66.74 71.335 67.5 ;
    RECT 71.815 66.74 72.035 67.5 ;
    RECT 72.515 66.74 72.735 67.5 ;
    RECT 73.215 66.74 73.435 67.5 ;
    RECT 73.915 66.74 74.835 67.5 ;
    RECT 75.315 66.74 75.535 67.5 ;
    RECT 76.015 66.74 76.225 67.5 ;
    RECT 76.705 66.74 76.92 67.5 ;
    RECT 77.4 66.74 77.62 67.5 ;
    RECT 78.1 66.74 78.32 67.5 ;
    RECT 78.8 66.74 79.02 67.5 ;
    RECT 79.5 66.74 81.115 67.5 ;
    RECT 81.595 66.74 81.815 67.5 ;
    RECT 82.295 66.74 82.515 67.5 ;
    RECT 82.995 66.74 83.055 67.5 ;
    RECT 83.055 66.65 83.335 67.59 ;
    RECT 83.335 66.74 83.505 67.5 ;
    RECT 26.71 65.98 26.88 66.74 ;
    RECT 26.88 65.89 27.16 66.83 ;
    RECT 27.16 65.98 27.32 66.74 ;
    RECT 27.8 65.98 28.02 66.74 ;
    RECT 28.5 65.98 28.72 66.74 ;
    RECT 29.2 65.98 30.815 66.74 ;
    RECT 31.295 65.98 31.515 66.74 ;
    RECT 31.995 65.98 32.21 66.74 ;
    RECT 32.69 65.98 32.91 66.74 ;
    RECT 33.39 65.98 33.61 66.74 ;
    RECT 34.09 65.98 34.31 66.74 ;
    RECT 34.79 65.98 35.005 66.74 ;
    RECT 35.485 65.98 36.405 66.74 ;
    RECT 36.885 65.98 37.105 66.74 ;
    RECT 37.585 65.98 37.8 66.74 ;
    RECT 38.28 65.98 38.5 66.74 ;
    RECT 38.98 65.98 39.2 66.74 ;
    RECT 39.68 65.98 39.895 66.74 ;
    RECT 40.375 65.98 40.595 66.74 ;
    RECT 41.075 65.98 41.995 66.74 ;
    RECT 42.475 65.98 42.69 66.74 ;
    RECT 43.17 65.98 43.39 66.74 ;
    RECT 43.87 65.98 44.09 66.74 ;
    RECT 44.57 65.98 44.79 66.74 ;
    RECT 45.27 65.98 45.485 66.74 ;
    RECT 45.965 65.98 46.185 66.74 ;
    RECT 46.665 65.98 47.58 66.74 ;
    RECT 48.06 65.98 48.28 66.74 ;
    RECT 48.76 65.98 48.98 66.74 ;
    RECT 49.46 65.98 49.68 66.74 ;
    RECT 50.16 65.98 50.375 66.74 ;
    RECT 50.855 65.98 51.775 66.74 ;
    RECT 52.255 65.98 53.17 66.74 ;
    RECT 53.65 65.98 53.87 66.74 ;
    RECT 54.35 65.98 54.57 66.74 ;
    RECT 55.05 65.98 55.265 66.74 ;
    RECT 55.745 65.98 55.965 66.74 ;
    RECT 56.445 65.98 56.665 66.74 ;
    RECT 57.145 65.98 58.06 66.74 ;
    RECT 58.54 65.98 59.46 66.74 ;
    RECT 59.94 65.98 60.16 66.74 ;
    RECT 60.64 65.98 60.855 66.74 ;
    RECT 61.335 65.98 61.555 66.74 ;
    RECT 62.035 65.98 62.25 66.74 ;
    RECT 62.73 65.98 63.65 66.74 ;
    RECT 64.13 65.98 64.345 66.74 ;
    RECT 64.825 65.98 65.045 66.74 ;
    RECT 65.525 65.98 65.745 66.74 ;
    RECT 66.225 65.98 66.445 66.74 ;
    RECT 66.925 65.98 67.14 66.74 ;
    RECT 67.62 65.98 67.84 66.74 ;
    RECT 68.32 65.98 69.235 66.74 ;
    RECT 69.715 65.98 69.935 66.74 ;
    RECT 70.415 65.98 70.635 66.74 ;
    RECT 71.115 65.98 71.335 66.74 ;
    RECT 71.815 65.98 72.035 66.74 ;
    RECT 72.515 65.98 72.735 66.74 ;
    RECT 73.215 65.98 73.435 66.74 ;
    RECT 73.915 65.98 74.835 66.74 ;
    RECT 75.315 65.98 75.535 66.74 ;
    RECT 76.015 65.98 76.225 66.74 ;
    RECT 76.705 65.98 76.92 66.74 ;
    RECT 77.4 65.98 77.62 66.74 ;
    RECT 78.1 65.98 78.32 66.74 ;
    RECT 78.8 65.98 79.02 66.74 ;
    RECT 79.5 65.98 81.115 66.74 ;
    RECT 81.595 65.98 81.815 66.74 ;
    RECT 82.295 65.98 82.515 66.74 ;
    RECT 82.995 65.98 83.055 66.74 ;
    RECT 83.055 65.89 83.335 66.83 ;
    RECT 83.335 65.98 83.505 66.74 ;
    RECT 26.71 65.22 26.88 65.98 ;
    RECT 26.88 65.13 27.16 66.07 ;
    RECT 27.16 65.22 27.32 65.98 ;
    RECT 27.8 65.22 28.02 65.98 ;
    RECT 28.5 65.22 28.72 65.98 ;
    RECT 29.2 65.22 30.815 65.98 ;
    RECT 31.295 65.22 31.515 65.98 ;
    RECT 31.995 65.22 32.21 65.98 ;
    RECT 32.69 65.22 32.91 65.98 ;
    RECT 33.39 65.22 33.61 65.98 ;
    RECT 34.09 65.22 34.31 65.98 ;
    RECT 34.79 65.22 35.005 65.98 ;
    RECT 35.485 65.22 36.405 65.98 ;
    RECT 36.885 65.22 37.105 65.98 ;
    RECT 37.585 65.22 37.8 65.98 ;
    RECT 38.28 65.22 38.5 65.98 ;
    RECT 38.98 65.22 39.2 65.98 ;
    RECT 39.68 65.22 39.895 65.98 ;
    RECT 40.375 65.22 40.595 65.98 ;
    RECT 41.075 65.22 41.995 65.98 ;
    RECT 42.475 65.22 42.69 65.98 ;
    RECT 43.17 65.22 43.39 65.98 ;
    RECT 43.87 65.22 44.09 65.98 ;
    RECT 44.57 65.22 44.79 65.98 ;
    RECT 45.27 65.22 45.485 65.98 ;
    RECT 45.965 65.22 46.185 65.98 ;
    RECT 46.665 65.22 47.58 65.98 ;
    RECT 48.06 65.22 48.28 65.98 ;
    RECT 48.76 65.22 48.98 65.98 ;
    RECT 49.46 65.22 49.68 65.98 ;
    RECT 50.16 65.22 50.375 65.98 ;
    RECT 50.855 65.22 51.775 65.98 ;
    RECT 52.255 65.22 53.17 65.98 ;
    RECT 53.65 65.22 53.87 65.98 ;
    RECT 54.35 65.22 54.57 65.98 ;
    RECT 55.05 65.22 55.265 65.98 ;
    RECT 55.745 65.22 55.965 65.98 ;
    RECT 56.445 65.22 56.665 65.98 ;
    RECT 57.145 65.22 58.06 65.98 ;
    RECT 58.54 65.22 59.46 65.98 ;
    RECT 59.94 65.22 60.16 65.98 ;
    RECT 60.64 65.22 60.855 65.98 ;
    RECT 61.335 65.22 61.555 65.98 ;
    RECT 62.035 65.22 62.25 65.98 ;
    RECT 62.73 65.22 63.65 65.98 ;
    RECT 64.13 65.22 64.345 65.98 ;
    RECT 64.825 65.22 65.045 65.98 ;
    RECT 65.525 65.22 65.745 65.98 ;
    RECT 66.225 65.22 66.445 65.98 ;
    RECT 66.925 65.22 67.14 65.98 ;
    RECT 67.62 65.22 67.84 65.98 ;
    RECT 68.32 65.22 69.235 65.98 ;
    RECT 69.715 65.22 69.935 65.98 ;
    RECT 70.415 65.22 70.635 65.98 ;
    RECT 71.115 65.22 71.335 65.98 ;
    RECT 71.815 65.22 72.035 65.98 ;
    RECT 72.515 65.22 72.735 65.98 ;
    RECT 73.215 65.22 73.435 65.98 ;
    RECT 73.915 65.22 74.835 65.98 ;
    RECT 75.315 65.22 75.535 65.98 ;
    RECT 76.015 65.22 76.225 65.98 ;
    RECT 76.705 65.22 76.92 65.98 ;
    RECT 77.4 65.22 77.62 65.98 ;
    RECT 78.1 65.22 78.32 65.98 ;
    RECT 78.8 65.22 79.02 65.98 ;
    RECT 79.5 65.22 81.115 65.98 ;
    RECT 81.595 65.22 81.815 65.98 ;
    RECT 82.295 65.22 82.515 65.98 ;
    RECT 82.995 65.22 83.055 65.98 ;
    RECT 83.055 65.13 83.335 66.07 ;
    RECT 83.335 65.22 83.505 65.98 ;
    RECT 26.71 64.46 26.88 65.22 ;
    RECT 26.88 64.37 27.16 65.31 ;
    RECT 27.16 64.46 27.32 65.22 ;
    RECT 27.8 64.46 28.02 65.22 ;
    RECT 28.5 64.46 28.72 65.22 ;
    RECT 29.2 64.46 30.815 65.22 ;
    RECT 31.295 64.46 31.515 65.22 ;
    RECT 31.995 64.46 32.21 65.22 ;
    RECT 32.69 64.46 32.91 65.22 ;
    RECT 33.39 64.46 33.61 65.22 ;
    RECT 34.09 64.46 34.31 65.22 ;
    RECT 34.79 64.46 35.005 65.22 ;
    RECT 35.485 64.46 36.405 65.22 ;
    RECT 36.885 64.46 37.105 65.22 ;
    RECT 37.585 64.46 37.8 65.22 ;
    RECT 38.28 64.46 38.5 65.22 ;
    RECT 38.98 64.46 39.2 65.22 ;
    RECT 39.68 64.46 39.895 65.22 ;
    RECT 40.375 64.46 40.595 65.22 ;
    RECT 41.075 64.46 41.995 65.22 ;
    RECT 42.475 64.46 42.69 65.22 ;
    RECT 43.17 64.46 43.39 65.22 ;
    RECT 43.87 64.46 44.09 65.22 ;
    RECT 44.57 64.46 44.79 65.22 ;
    RECT 45.27 64.46 45.485 65.22 ;
    RECT 45.965 64.46 46.185 65.22 ;
    RECT 46.665 64.46 47.58 65.22 ;
    RECT 48.06 64.46 48.28 65.22 ;
    RECT 48.76 64.46 48.98 65.22 ;
    RECT 49.46 64.46 49.68 65.22 ;
    RECT 50.16 64.46 50.375 65.22 ;
    RECT 50.855 64.46 51.775 65.22 ;
    RECT 52.255 64.46 53.17 65.22 ;
    RECT 53.65 64.46 53.87 65.22 ;
    RECT 54.35 64.46 54.57 65.22 ;
    RECT 55.05 64.46 55.265 65.22 ;
    RECT 55.745 64.46 55.965 65.22 ;
    RECT 56.445 64.46 56.665 65.22 ;
    RECT 57.145 64.46 58.06 65.22 ;
    RECT 58.54 64.46 59.46 65.22 ;
    RECT 59.94 64.46 60.16 65.22 ;
    RECT 60.64 64.46 60.855 65.22 ;
    RECT 61.335 64.46 61.555 65.22 ;
    RECT 62.035 64.46 62.25 65.22 ;
    RECT 62.73 64.46 63.65 65.22 ;
    RECT 64.13 64.46 64.345 65.22 ;
    RECT 64.825 64.46 65.045 65.22 ;
    RECT 65.525 64.46 65.745 65.22 ;
    RECT 66.225 64.46 66.445 65.22 ;
    RECT 66.925 64.46 67.14 65.22 ;
    RECT 67.62 64.46 67.84 65.22 ;
    RECT 68.32 64.46 69.235 65.22 ;
    RECT 69.715 64.46 69.935 65.22 ;
    RECT 70.415 64.46 70.635 65.22 ;
    RECT 71.115 64.46 71.335 65.22 ;
    RECT 71.815 64.46 72.035 65.22 ;
    RECT 72.515 64.46 72.735 65.22 ;
    RECT 73.215 64.46 73.435 65.22 ;
    RECT 73.915 64.46 74.835 65.22 ;
    RECT 75.315 64.46 75.535 65.22 ;
    RECT 76.015 64.46 76.225 65.22 ;
    RECT 76.705 64.46 76.92 65.22 ;
    RECT 77.4 64.46 77.62 65.22 ;
    RECT 78.1 64.46 78.32 65.22 ;
    RECT 78.8 64.46 79.02 65.22 ;
    RECT 79.5 64.46 81.115 65.22 ;
    RECT 81.595 64.46 81.815 65.22 ;
    RECT 82.295 64.46 82.515 65.22 ;
    RECT 82.995 64.46 83.055 65.22 ;
    RECT 83.055 64.37 83.335 65.31 ;
    RECT 83.335 64.46 83.505 65.22 ;
    RECT 26.71 63.7 26.88 64.46 ;
    RECT 26.88 63.61 27.16 64.55 ;
    RECT 27.16 63.7 27.32 64.46 ;
    RECT 27.8 63.7 28.02 64.46 ;
    RECT 28.5 63.7 28.72 64.46 ;
    RECT 29.2 63.7 30.815 64.46 ;
    RECT 31.295 63.7 31.515 64.46 ;
    RECT 31.995 63.7 32.21 64.46 ;
    RECT 32.69 63.7 32.91 64.46 ;
    RECT 33.39 63.7 33.61 64.46 ;
    RECT 34.09 63.7 34.31 64.46 ;
    RECT 34.79 63.7 35.005 64.46 ;
    RECT 35.485 63.7 36.405 64.46 ;
    RECT 36.885 63.7 37.105 64.46 ;
    RECT 37.585 63.7 37.8 64.46 ;
    RECT 38.28 63.7 38.5 64.46 ;
    RECT 38.98 63.7 39.2 64.46 ;
    RECT 39.68 63.7 39.895 64.46 ;
    RECT 40.375 63.7 40.595 64.46 ;
    RECT 41.075 63.7 41.995 64.46 ;
    RECT 42.475 63.7 42.69 64.46 ;
    RECT 43.17 63.7 43.39 64.46 ;
    RECT 43.87 63.7 44.09 64.46 ;
    RECT 44.57 63.7 44.79 64.46 ;
    RECT 45.27 63.7 45.485 64.46 ;
    RECT 45.965 63.7 46.185 64.46 ;
    RECT 46.665 63.7 47.58 64.46 ;
    RECT 48.06 63.7 48.28 64.46 ;
    RECT 48.76 63.7 48.98 64.46 ;
    RECT 49.46 63.7 49.68 64.46 ;
    RECT 50.16 63.7 50.375 64.46 ;
    RECT 50.855 63.7 51.775 64.46 ;
    RECT 52.255 63.7 53.17 64.46 ;
    RECT 53.65 63.7 53.87 64.46 ;
    RECT 54.35 63.7 54.57 64.46 ;
    RECT 55.05 63.7 55.265 64.46 ;
    RECT 55.745 63.7 55.965 64.46 ;
    RECT 56.445 63.7 56.665 64.46 ;
    RECT 57.145 63.7 58.06 64.46 ;
    RECT 58.54 63.7 59.46 64.46 ;
    RECT 59.94 63.7 60.16 64.46 ;
    RECT 60.64 63.7 60.855 64.46 ;
    RECT 61.335 63.7 61.555 64.46 ;
    RECT 62.035 63.7 62.25 64.46 ;
    RECT 62.73 63.7 63.65 64.46 ;
    RECT 64.13 63.7 64.345 64.46 ;
    RECT 64.825 63.7 65.045 64.46 ;
    RECT 65.525 63.7 65.745 64.46 ;
    RECT 66.225 63.7 66.445 64.46 ;
    RECT 66.925 63.7 67.14 64.46 ;
    RECT 67.62 63.7 67.84 64.46 ;
    RECT 68.32 63.7 69.235 64.46 ;
    RECT 69.715 63.7 69.935 64.46 ;
    RECT 70.415 63.7 70.635 64.46 ;
    RECT 71.115 63.7 71.335 64.46 ;
    RECT 71.815 63.7 72.035 64.46 ;
    RECT 72.515 63.7 72.735 64.46 ;
    RECT 73.215 63.7 73.435 64.46 ;
    RECT 73.915 63.7 74.835 64.46 ;
    RECT 75.315 63.7 75.535 64.46 ;
    RECT 76.015 63.7 76.225 64.46 ;
    RECT 76.705 63.7 76.92 64.46 ;
    RECT 77.4 63.7 77.62 64.46 ;
    RECT 78.1 63.7 78.32 64.46 ;
    RECT 78.8 63.7 79.02 64.46 ;
    RECT 79.5 63.7 81.115 64.46 ;
    RECT 81.595 63.7 81.815 64.46 ;
    RECT 82.295 63.7 82.515 64.46 ;
    RECT 82.995 63.7 83.055 64.46 ;
    RECT 83.055 63.61 83.335 64.55 ;
    RECT 83.335 63.7 83.505 64.46 ;
    RECT 26.71 62.94 26.88 63.7 ;
    RECT 26.88 62.85 27.16 63.79 ;
    RECT 27.16 62.94 27.32 63.7 ;
    RECT 27.8 62.94 28.02 63.7 ;
    RECT 28.5 62.94 28.72 63.7 ;
    RECT 29.2 62.94 30.815 63.7 ;
    RECT 31.295 62.94 31.515 63.7 ;
    RECT 31.995 62.94 32.21 63.7 ;
    RECT 32.69 62.94 32.91 63.7 ;
    RECT 33.39 62.94 33.61 63.7 ;
    RECT 34.09 62.94 34.31 63.7 ;
    RECT 34.79 62.94 35.005 63.7 ;
    RECT 35.485 62.94 36.405 63.7 ;
    RECT 36.885 62.94 37.105 63.7 ;
    RECT 37.585 62.94 37.8 63.7 ;
    RECT 38.28 62.94 38.5 63.7 ;
    RECT 38.98 62.94 39.2 63.7 ;
    RECT 39.68 62.94 39.895 63.7 ;
    RECT 40.375 62.94 40.595 63.7 ;
    RECT 41.075 62.94 41.995 63.7 ;
    RECT 42.475 62.94 42.69 63.7 ;
    RECT 43.17 62.94 43.39 63.7 ;
    RECT 43.87 62.94 44.09 63.7 ;
    RECT 44.57 62.94 44.79 63.7 ;
    RECT 45.27 62.94 45.485 63.7 ;
    RECT 45.965 62.94 46.185 63.7 ;
    RECT 46.665 62.94 47.58 63.7 ;
    RECT 48.06 62.94 48.28 63.7 ;
    RECT 48.76 62.94 48.98 63.7 ;
    RECT 49.46 62.94 49.68 63.7 ;
    RECT 50.16 62.94 50.375 63.7 ;
    RECT 50.855 62.94 51.775 63.7 ;
    RECT 52.255 62.94 53.17 63.7 ;
    RECT 53.65 62.94 53.87 63.7 ;
    RECT 54.35 62.94 54.57 63.7 ;
    RECT 55.05 62.94 55.265 63.7 ;
    RECT 55.745 62.94 55.965 63.7 ;
    RECT 56.445 62.94 56.665 63.7 ;
    RECT 57.145 62.94 58.06 63.7 ;
    RECT 58.54 62.94 59.46 63.7 ;
    RECT 59.94 62.94 60.16 63.7 ;
    RECT 60.64 62.94 60.855 63.7 ;
    RECT 61.335 62.94 61.555 63.7 ;
    RECT 62.035 62.94 62.25 63.7 ;
    RECT 62.73 62.94 63.65 63.7 ;
    RECT 64.13 62.94 64.345 63.7 ;
    RECT 64.825 62.94 65.045 63.7 ;
    RECT 65.525 62.94 65.745 63.7 ;
    RECT 66.225 62.94 66.445 63.7 ;
    RECT 66.925 62.94 67.14 63.7 ;
    RECT 67.62 62.94 67.84 63.7 ;
    RECT 68.32 62.94 69.235 63.7 ;
    RECT 69.715 62.94 69.935 63.7 ;
    RECT 70.415 62.94 70.635 63.7 ;
    RECT 71.115 62.94 71.335 63.7 ;
    RECT 71.815 62.94 72.035 63.7 ;
    RECT 72.515 62.94 72.735 63.7 ;
    RECT 73.215 62.94 73.435 63.7 ;
    RECT 73.915 62.94 74.835 63.7 ;
    RECT 75.315 62.94 75.535 63.7 ;
    RECT 76.015 62.94 76.225 63.7 ;
    RECT 76.705 62.94 76.92 63.7 ;
    RECT 77.4 62.94 77.62 63.7 ;
    RECT 78.1 62.94 78.32 63.7 ;
    RECT 78.8 62.94 79.02 63.7 ;
    RECT 79.5 62.94 81.115 63.7 ;
    RECT 81.595 62.94 81.815 63.7 ;
    RECT 82.295 62.94 82.515 63.7 ;
    RECT 82.995 62.94 83.055 63.7 ;
    RECT 83.055 62.85 83.335 63.79 ;
    RECT 83.335 62.94 83.505 63.7 ;
    RECT 26.71 62.18 26.88 62.94 ;
    RECT 26.88 62.09 27.16 63.03 ;
    RECT 27.16 62.18 27.32 62.94 ;
    RECT 27.8 62.18 28.02 62.94 ;
    RECT 28.5 62.18 28.72 62.94 ;
    RECT 29.2 62.18 30.815 62.94 ;
    RECT 31.295 62.18 31.515 62.94 ;
    RECT 31.995 62.18 32.21 62.94 ;
    RECT 32.69 62.18 32.91 62.94 ;
    RECT 33.39 62.18 33.61 62.94 ;
    RECT 34.09 62.18 34.31 62.94 ;
    RECT 34.79 62.18 35.005 62.94 ;
    RECT 35.485 62.18 36.405 62.94 ;
    RECT 36.885 62.18 37.105 62.94 ;
    RECT 37.585 62.18 37.8 62.94 ;
    RECT 38.28 62.18 38.5 62.94 ;
    RECT 38.98 62.18 39.2 62.94 ;
    RECT 39.68 62.18 39.895 62.94 ;
    RECT 40.375 62.18 40.595 62.94 ;
    RECT 41.075 62.18 41.995 62.94 ;
    RECT 42.475 62.18 42.69 62.94 ;
    RECT 43.17 62.18 43.39 62.94 ;
    RECT 43.87 62.18 44.09 62.94 ;
    RECT 44.57 62.18 44.79 62.94 ;
    RECT 45.27 62.18 45.485 62.94 ;
    RECT 45.965 62.18 46.185 62.94 ;
    RECT 46.665 62.18 47.58 62.94 ;
    RECT 48.06 62.18 48.28 62.94 ;
    RECT 48.76 62.18 48.98 62.94 ;
    RECT 49.46 62.18 49.68 62.94 ;
    RECT 50.16 62.18 50.375 62.94 ;
    RECT 50.855 62.18 51.775 62.94 ;
    RECT 52.255 62.18 53.17 62.94 ;
    RECT 53.65 62.18 53.87 62.94 ;
    RECT 54.35 62.18 54.57 62.94 ;
    RECT 55.05 62.18 55.265 62.94 ;
    RECT 55.745 62.18 55.965 62.94 ;
    RECT 56.445 62.18 56.665 62.94 ;
    RECT 57.145 62.18 58.06 62.94 ;
    RECT 58.54 62.18 59.46 62.94 ;
    RECT 59.94 62.18 60.16 62.94 ;
    RECT 60.64 62.18 60.855 62.94 ;
    RECT 61.335 62.18 61.555 62.94 ;
    RECT 62.035 62.18 62.25 62.94 ;
    RECT 62.73 62.18 63.65 62.94 ;
    RECT 64.13 62.18 64.345 62.94 ;
    RECT 64.825 62.18 65.045 62.94 ;
    RECT 65.525 62.18 65.745 62.94 ;
    RECT 66.225 62.18 66.445 62.94 ;
    RECT 66.925 62.18 67.14 62.94 ;
    RECT 67.62 62.18 67.84 62.94 ;
    RECT 68.32 62.18 69.235 62.94 ;
    RECT 69.715 62.18 69.935 62.94 ;
    RECT 70.415 62.18 70.635 62.94 ;
    RECT 71.115 62.18 71.335 62.94 ;
    RECT 71.815 62.18 72.035 62.94 ;
    RECT 72.515 62.18 72.735 62.94 ;
    RECT 73.215 62.18 73.435 62.94 ;
    RECT 73.915 62.18 74.835 62.94 ;
    RECT 75.315 62.18 75.535 62.94 ;
    RECT 76.015 62.18 76.225 62.94 ;
    RECT 76.705 62.18 76.92 62.94 ;
    RECT 77.4 62.18 77.62 62.94 ;
    RECT 78.1 62.18 78.32 62.94 ;
    RECT 78.8 62.18 79.02 62.94 ;
    RECT 79.5 62.18 81.115 62.94 ;
    RECT 81.595 62.18 81.815 62.94 ;
    RECT 82.295 62.18 82.515 62.94 ;
    RECT 82.995 62.18 83.055 62.94 ;
    RECT 83.055 62.09 83.335 63.03 ;
    RECT 83.335 62.18 83.505 62.94 ;
    RECT 26.71 61.42 26.88 62.18 ;
    RECT 26.88 61.33 27.16 62.27 ;
    RECT 27.16 61.42 27.32 62.18 ;
    RECT 27.8 61.42 28.02 62.18 ;
    RECT 28.5 61.42 28.72 62.18 ;
    RECT 29.2 61.42 30.815 62.18 ;
    RECT 31.295 61.42 31.515 62.18 ;
    RECT 31.995 61.42 32.21 62.18 ;
    RECT 32.69 61.42 32.91 62.18 ;
    RECT 33.39 61.42 33.61 62.18 ;
    RECT 34.09 61.42 34.31 62.18 ;
    RECT 34.79 61.42 35.005 62.18 ;
    RECT 35.485 61.42 36.405 62.18 ;
    RECT 36.885 61.42 37.105 62.18 ;
    RECT 37.585 61.42 37.8 62.18 ;
    RECT 38.28 61.42 38.5 62.18 ;
    RECT 38.98 61.42 39.2 62.18 ;
    RECT 39.68 61.42 39.895 62.18 ;
    RECT 40.375 61.42 40.595 62.18 ;
    RECT 41.075 61.42 41.995 62.18 ;
    RECT 42.475 61.42 42.69 62.18 ;
    RECT 43.17 61.42 43.39 62.18 ;
    RECT 43.87 61.42 44.09 62.18 ;
    RECT 44.57 61.42 44.79 62.18 ;
    RECT 45.27 61.42 45.485 62.18 ;
    RECT 45.965 61.42 46.185 62.18 ;
    RECT 46.665 61.42 47.58 62.18 ;
    RECT 48.06 61.42 48.28 62.18 ;
    RECT 48.76 61.42 48.98 62.18 ;
    RECT 49.46 61.42 49.68 62.18 ;
    RECT 50.16 61.42 50.375 62.18 ;
    RECT 50.855 61.42 51.775 62.18 ;
    RECT 52.255 61.42 53.17 62.18 ;
    RECT 53.65 61.42 53.87 62.18 ;
    RECT 54.35 61.42 54.57 62.18 ;
    RECT 55.05 61.42 55.265 62.18 ;
    RECT 55.745 61.42 55.965 62.18 ;
    RECT 56.445 61.42 56.665 62.18 ;
    RECT 57.145 61.42 58.06 62.18 ;
    RECT 58.54 61.42 59.46 62.18 ;
    RECT 59.94 61.42 60.16 62.18 ;
    RECT 60.64 61.42 60.855 62.18 ;
    RECT 61.335 61.42 61.555 62.18 ;
    RECT 62.035 61.42 62.25 62.18 ;
    RECT 62.73 61.42 63.65 62.18 ;
    RECT 64.13 61.42 64.345 62.18 ;
    RECT 64.825 61.42 65.045 62.18 ;
    RECT 65.525 61.42 65.745 62.18 ;
    RECT 66.225 61.42 66.445 62.18 ;
    RECT 66.925 61.42 67.14 62.18 ;
    RECT 67.62 61.42 67.84 62.18 ;
    RECT 68.32 61.42 69.235 62.18 ;
    RECT 69.715 61.42 69.935 62.18 ;
    RECT 70.415 61.42 70.635 62.18 ;
    RECT 71.115 61.42 71.335 62.18 ;
    RECT 71.815 61.42 72.035 62.18 ;
    RECT 72.515 61.42 72.735 62.18 ;
    RECT 73.215 61.42 73.435 62.18 ;
    RECT 73.915 61.42 74.835 62.18 ;
    RECT 75.315 61.42 75.535 62.18 ;
    RECT 76.015 61.42 76.225 62.18 ;
    RECT 76.705 61.42 76.92 62.18 ;
    RECT 77.4 61.42 77.62 62.18 ;
    RECT 78.1 61.42 78.32 62.18 ;
    RECT 78.8 61.42 79.02 62.18 ;
    RECT 79.5 61.42 81.115 62.18 ;
    RECT 81.595 61.42 81.815 62.18 ;
    RECT 82.295 61.42 82.515 62.18 ;
    RECT 82.995 61.42 83.055 62.18 ;
    RECT 83.055 61.33 83.335 62.27 ;
    RECT 83.335 61.42 83.505 62.18 ;
    RECT 26.71 60.66 26.88 61.42 ;
    RECT 26.88 60.57 27.16 61.51 ;
    RECT 27.16 60.66 27.32 61.42 ;
    RECT 27.8 60.66 28.02 61.42 ;
    RECT 28.5 60.66 28.72 61.42 ;
    RECT 29.2 60.66 30.815 61.42 ;
    RECT 31.295 60.66 31.515 61.42 ;
    RECT 31.995 60.66 32.21 61.42 ;
    RECT 32.69 60.66 32.91 61.42 ;
    RECT 33.39 60.66 33.61 61.42 ;
    RECT 34.09 60.66 34.31 61.42 ;
    RECT 34.79 60.66 35.005 61.42 ;
    RECT 35.485 60.66 36.405 61.42 ;
    RECT 36.885 60.66 37.105 61.42 ;
    RECT 37.585 60.66 37.8 61.42 ;
    RECT 38.28 60.66 38.5 61.42 ;
    RECT 38.98 60.66 39.2 61.42 ;
    RECT 39.68 60.66 39.895 61.42 ;
    RECT 40.375 60.66 40.595 61.42 ;
    RECT 41.075 60.66 41.995 61.42 ;
    RECT 42.475 60.66 42.69 61.42 ;
    RECT 43.17 60.66 43.39 61.42 ;
    RECT 43.87 60.66 44.09 61.42 ;
    RECT 44.57 60.66 44.79 61.42 ;
    RECT 45.27 60.66 45.485 61.42 ;
    RECT 45.965 60.66 46.185 61.42 ;
    RECT 46.665 60.66 47.58 61.42 ;
    RECT 48.06 60.66 48.28 61.42 ;
    RECT 48.76 60.66 48.98 61.42 ;
    RECT 49.46 60.66 49.68 61.42 ;
    RECT 50.16 60.66 50.375 61.42 ;
    RECT 50.855 60.66 51.775 61.42 ;
    RECT 52.255 60.66 53.17 61.42 ;
    RECT 53.65 60.66 53.87 61.42 ;
    RECT 54.35 60.66 54.57 61.42 ;
    RECT 55.05 60.66 55.265 61.42 ;
    RECT 55.745 60.66 55.965 61.42 ;
    RECT 56.445 60.66 56.665 61.42 ;
    RECT 57.145 60.66 58.06 61.42 ;
    RECT 58.54 60.66 59.46 61.42 ;
    RECT 59.94 60.66 60.16 61.42 ;
    RECT 60.64 60.66 60.855 61.42 ;
    RECT 61.335 60.66 61.555 61.42 ;
    RECT 62.035 60.66 62.25 61.42 ;
    RECT 62.73 60.66 63.65 61.42 ;
    RECT 64.13 60.66 64.345 61.42 ;
    RECT 64.825 60.66 65.045 61.42 ;
    RECT 65.525 60.66 65.745 61.42 ;
    RECT 66.225 60.66 66.445 61.42 ;
    RECT 66.925 60.66 67.14 61.42 ;
    RECT 67.62 60.66 67.84 61.42 ;
    RECT 68.32 60.66 69.235 61.42 ;
    RECT 69.715 60.66 69.935 61.42 ;
    RECT 70.415 60.66 70.635 61.42 ;
    RECT 71.115 60.66 71.335 61.42 ;
    RECT 71.815 60.66 72.035 61.42 ;
    RECT 72.515 60.66 72.735 61.42 ;
    RECT 73.215 60.66 73.435 61.42 ;
    RECT 73.915 60.66 74.835 61.42 ;
    RECT 75.315 60.66 75.535 61.42 ;
    RECT 76.015 60.66 76.225 61.42 ;
    RECT 76.705 60.66 76.92 61.42 ;
    RECT 77.4 60.66 77.62 61.42 ;
    RECT 78.1 60.66 78.32 61.42 ;
    RECT 78.8 60.66 79.02 61.42 ;
    RECT 79.5 60.66 81.115 61.42 ;
    RECT 81.595 60.66 81.815 61.42 ;
    RECT 82.295 60.66 82.515 61.42 ;
    RECT 82.995 60.66 83.055 61.42 ;
    RECT 83.055 60.57 83.335 61.51 ;
    RECT 83.335 60.66 83.505 61.42 ;
    RECT 26.71 59.92 26.88 60.66 ;
    RECT 26.88 59.785 27.16 60.81 ;
    RECT 27.16 59.92 27.32 60.66 ;
    RECT 27.8 59.92 28.02 60.66 ;
    RECT 28.5 59.92 28.72 60.66 ;
    RECT 29.2 59.92 29.52 60.66 ;
    RECT 29.52 59.86 29.8 60.725 ;
    RECT 29.8 59.92 30.215 60.66 ;
    RECT 30.215 59.86 30.495 60.725 ;
    RECT 30.495 59.92 30.615 60.66 ;
    RECT 30.615 59.86 30.795 60.725 ;
    RECT 30.795 59.92 30.815 60.66 ;
    RECT 31.295 59.92 31.515 60.66 ;
    RECT 31.995 59.92 32.21 60.66 ;
    RECT 32.69 59.92 32.91 60.66 ;
    RECT 33.39 59.92 33.61 60.66 ;
    RECT 34.09 59.92 34.31 60.66 ;
    RECT 34.79 59.92 35.005 60.66 ;
    RECT 35.485 59.92 35.805 60.66 ;
    RECT 35.805 59.86 36.085 60.725 ;
    RECT 36.085 59.92 36.405 60.66 ;
    RECT 36.885 59.92 37.105 60.66 ;
    RECT 37.585 59.92 37.8 60.66 ;
    RECT 38.28 59.92 38.5 60.66 ;
    RECT 38.98 59.92 39.2 60.66 ;
    RECT 39.68 59.92 39.895 60.66 ;
    RECT 40.375 59.92 40.595 60.66 ;
    RECT 41.075 59.92 41.395 60.66 ;
    RECT 41.395 59.86 41.675 60.725 ;
    RECT 41.675 59.92 41.995 60.66 ;
    RECT 42.475 59.92 42.69 60.66 ;
    RECT 43.17 59.92 43.39 60.66 ;
    RECT 43.87 59.92 44.09 60.66 ;
    RECT 44.57 59.92 44.79 60.66 ;
    RECT 45.27 59.92 45.485 60.66 ;
    RECT 45.965 59.92 46.185 60.66 ;
    RECT 46.665 59.92 46.985 60.66 ;
    RECT 46.985 59.86 47.265 60.725 ;
    RECT 47.265 59.92 47.58 60.66 ;
    RECT 48.06 59.92 48.28 60.66 ;
    RECT 48.76 59.92 48.98 60.66 ;
    RECT 49.46 59.92 49.68 60.66 ;
    RECT 50.16 59.92 50.375 60.66 ;
    RECT 50.855 59.92 50.875 60.66 ;
    RECT 50.875 59.86 51.055 60.725 ;
    RECT 51.055 59.92 51.175 60.66 ;
    RECT 51.175 59.86 51.455 60.725 ;
    RECT 51.455 59.92 51.775 60.66 ;
    RECT 52.255 59.92 52.575 60.66 ;
    RECT 52.575 59.86 52.855 60.725 ;
    RECT 52.855 59.92 53.17 60.66 ;
    RECT 53.65 59.92 53.87 60.66 ;
    RECT 54.35 59.92 54.57 60.66 ;
    RECT 55.05 59.92 55.265 60.66 ;
    RECT 55.745 59.92 55.965 60.66 ;
    RECT 56.445 59.92 56.665 60.66 ;
    RECT 57.145 59.92 57.465 60.66 ;
    RECT 57.465 59.86 57.745 60.725 ;
    RECT 57.745 59.92 58.06 60.66 ;
    RECT 58.54 59.92 58.86 60.66 ;
    RECT 58.86 59.86 59.14 60.725 ;
    RECT 59.14 59.92 59.26 60.66 ;
    RECT 59.26 59.86 59.44 60.725 ;
    RECT 59.44 59.92 59.46 60.66 ;
    RECT 59.94 59.92 60.16 60.66 ;
    RECT 60.64 59.92 60.855 60.66 ;
    RECT 61.335 59.92 61.555 60.66 ;
    RECT 62.035 59.92 62.25 60.66 ;
    RECT 62.73 59.92 63.05 60.66 ;
    RECT 63.05 59.86 63.33 60.725 ;
    RECT 63.33 59.92 63.65 60.66 ;
    RECT 64.13 59.92 64.345 60.66 ;
    RECT 64.825 59.92 65.045 60.66 ;
    RECT 65.525 59.92 65.745 60.66 ;
    RECT 66.225 59.92 66.445 60.66 ;
    RECT 66.925 59.92 67.14 60.66 ;
    RECT 67.62 59.92 67.84 60.66 ;
    RECT 68.32 59.92 68.64 60.66 ;
    RECT 68.64 59.86 68.92 60.725 ;
    RECT 68.92 59.92 69.235 60.66 ;
    RECT 69.715 59.92 69.935 60.66 ;
    RECT 70.415 59.92 70.635 60.66 ;
    RECT 71.115 59.92 71.335 60.66 ;
    RECT 71.815 59.92 72.035 60.66 ;
    RECT 72.515 59.92 72.735 60.66 ;
    RECT 73.215 59.92 73.435 60.66 ;
    RECT 73.915 59.92 74.235 60.66 ;
    RECT 74.235 59.86 74.515 60.725 ;
    RECT 74.515 59.92 74.835 60.66 ;
    RECT 75.315 59.92 75.535 60.66 ;
    RECT 76.015 59.92 76.07 60.66 ;
    RECT 76.07 59.86 76.17 60.725 ;
    RECT 76.17 59.92 76.225 60.66 ;
    RECT 76.705 59.92 76.765 60.66 ;
    RECT 76.765 59.86 76.865 60.725 ;
    RECT 76.865 59.92 76.92 60.66 ;
    RECT 77.4 59.92 77.62 60.66 ;
    RECT 78.1 59.92 78.32 60.66 ;
    RECT 78.8 59.92 79.02 60.66 ;
    RECT 79.5 59.92 79.52 60.66 ;
    RECT 79.52 59.86 79.7 60.725 ;
    RECT 79.7 59.92 79.82 60.66 ;
    RECT 79.82 59.86 80.1 60.725 ;
    RECT 80.1 59.92 80.515 60.66 ;
    RECT 80.515 59.86 80.795 60.725 ;
    RECT 80.795 59.92 81.115 60.66 ;
    RECT 81.595 59.92 81.815 60.66 ;
    RECT 82.295 59.92 82.515 60.66 ;
    RECT 82.995 59.92 83.055 60.66 ;
    RECT 83.055 59.77 83.335 60.81 ;
    RECT 83.335 59.92 83.505 60.66 ;
    RECT 26.71 59.16 26.88 59.92 ;
    RECT 26.88 59.07 27.16 60.01 ;
    RECT 27.16 59.16 27.32 59.92 ;
    RECT 27.8 59.16 28.02 59.92 ;
    RECT 28.5 59.16 28.72 59.92 ;
    RECT 29.2 59.16 30.815 59.92 ;
    RECT 31.295 59.16 31.515 59.92 ;
    RECT 31.995 59.16 32.21 59.92 ;
    RECT 32.69 59.16 32.91 59.92 ;
    RECT 33.39 59.16 33.61 59.92 ;
    RECT 34.09 59.16 34.31 59.92 ;
    RECT 34.79 59.16 35.005 59.92 ;
    RECT 35.485 59.16 36.405 59.92 ;
    RECT 36.885 59.16 37.105 59.92 ;
    RECT 37.585 59.16 37.8 59.92 ;
    RECT 38.28 59.16 38.5 59.92 ;
    RECT 38.98 59.16 39.2 59.92 ;
    RECT 39.68 59.16 39.895 59.92 ;
    RECT 40.375 59.16 40.595 59.92 ;
    RECT 41.075 59.16 41.995 59.92 ;
    RECT 42.475 59.16 42.69 59.92 ;
    RECT 43.17 59.16 43.39 59.92 ;
    RECT 43.87 59.16 44.09 59.92 ;
    RECT 44.57 59.16 44.79 59.92 ;
    RECT 45.27 59.16 45.485 59.92 ;
    RECT 45.965 59.16 46.185 59.92 ;
    RECT 46.665 59.16 47.58 59.92 ;
    RECT 48.06 59.16 48.28 59.92 ;
    RECT 48.76 59.16 48.98 59.92 ;
    RECT 49.46 59.16 49.68 59.92 ;
    RECT 50.16 59.16 50.375 59.92 ;
    RECT 50.855 59.16 51.775 59.92 ;
    RECT 52.255 59.16 53.17 59.92 ;
    RECT 53.65 59.16 53.87 59.92 ;
    RECT 54.35 59.16 54.57 59.92 ;
    RECT 55.05 59.16 55.265 59.92 ;
    RECT 55.745 59.16 55.965 59.92 ;
    RECT 56.445 59.16 56.665 59.92 ;
    RECT 57.145 59.16 58.06 59.92 ;
    RECT 58.54 59.16 59.46 59.92 ;
    RECT 59.94 59.16 60.16 59.92 ;
    RECT 60.64 59.16 60.855 59.92 ;
    RECT 61.335 59.16 61.555 59.92 ;
    RECT 62.035 59.16 62.25 59.92 ;
    RECT 62.73 59.16 63.65 59.92 ;
    RECT 64.13 59.16 64.345 59.92 ;
    RECT 64.825 59.16 65.045 59.92 ;
    RECT 65.525 59.16 65.745 59.92 ;
    RECT 66.225 59.16 66.445 59.92 ;
    RECT 66.925 59.16 67.14 59.92 ;
    RECT 67.62 59.16 67.84 59.92 ;
    RECT 68.32 59.16 69.235 59.92 ;
    RECT 69.715 59.16 69.935 59.92 ;
    RECT 70.415 59.16 70.635 59.92 ;
    RECT 71.115 59.16 71.335 59.92 ;
    RECT 71.815 59.16 72.035 59.92 ;
    RECT 72.515 59.16 72.735 59.92 ;
    RECT 73.215 59.16 73.435 59.92 ;
    RECT 73.915 59.16 74.835 59.92 ;
    RECT 75.315 59.16 75.535 59.92 ;
    RECT 76.015 59.16 76.225 59.92 ;
    RECT 76.705 59.16 76.92 59.92 ;
    RECT 77.4 59.16 77.62 59.92 ;
    RECT 78.1 59.16 78.32 59.92 ;
    RECT 78.8 59.16 79.02 59.92 ;
    RECT 79.5 59.16 81.115 59.92 ;
    RECT 81.595 59.16 81.815 59.92 ;
    RECT 82.295 59.16 82.515 59.92 ;
    RECT 82.995 59.16 83.055 59.92 ;
    RECT 83.055 59.07 83.335 60.01 ;
    RECT 83.335 59.16 83.505 59.92 ;
    RECT 26.71 58.4 26.88 59.16 ;
    RECT 26.88 58.31 27.16 59.25 ;
    RECT 27.16 58.4 27.32 59.16 ;
    RECT 27.8 58.4 28.02 59.16 ;
    RECT 28.5 58.4 28.72 59.16 ;
    RECT 29.2 58.4 30.815 59.16 ;
    RECT 31.295 58.4 31.515 59.16 ;
    RECT 31.995 58.4 32.21 59.16 ;
    RECT 32.69 58.4 32.91 59.16 ;
    RECT 33.39 58.4 33.61 59.16 ;
    RECT 34.09 58.4 34.31 59.16 ;
    RECT 34.79 58.4 35.005 59.16 ;
    RECT 35.485 58.4 36.405 59.16 ;
    RECT 36.885 58.4 37.105 59.16 ;
    RECT 37.585 58.4 37.8 59.16 ;
    RECT 38.28 58.4 38.5 59.16 ;
    RECT 38.98 58.4 39.2 59.16 ;
    RECT 39.68 58.4 39.895 59.16 ;
    RECT 40.375 58.4 40.595 59.16 ;
    RECT 41.075 58.4 41.995 59.16 ;
    RECT 42.475 58.4 42.69 59.16 ;
    RECT 43.17 58.4 43.39 59.16 ;
    RECT 43.87 58.4 44.09 59.16 ;
    RECT 44.57 58.4 44.79 59.16 ;
    RECT 45.27 58.4 45.485 59.16 ;
    RECT 45.965 58.4 46.185 59.16 ;
    RECT 46.665 58.4 47.58 59.16 ;
    RECT 48.06 58.4 48.28 59.16 ;
    RECT 48.76 58.4 48.98 59.16 ;
    RECT 49.46 58.4 49.68 59.16 ;
    RECT 50.16 58.4 50.375 59.16 ;
    RECT 50.855 58.4 51.775 59.16 ;
    RECT 52.255 58.4 53.17 59.16 ;
    RECT 53.65 58.4 53.87 59.16 ;
    RECT 54.35 58.4 54.57 59.16 ;
    RECT 55.05 58.4 55.265 59.16 ;
    RECT 55.745 58.4 55.965 59.16 ;
    RECT 56.445 58.4 56.665 59.16 ;
    RECT 57.145 58.4 58.06 59.16 ;
    RECT 58.54 58.4 59.46 59.16 ;
    RECT 59.94 58.4 60.16 59.16 ;
    RECT 60.64 58.4 60.855 59.16 ;
    RECT 61.335 58.4 61.555 59.16 ;
    RECT 62.035 58.4 62.25 59.16 ;
    RECT 62.73 58.4 63.65 59.16 ;
    RECT 64.13 58.4 64.345 59.16 ;
    RECT 64.825 58.4 65.045 59.16 ;
    RECT 65.525 58.4 65.745 59.16 ;
    RECT 66.225 58.4 66.445 59.16 ;
    RECT 66.925 58.4 67.14 59.16 ;
    RECT 67.62 58.4 67.84 59.16 ;
    RECT 68.32 58.4 69.235 59.16 ;
    RECT 69.715 58.4 69.935 59.16 ;
    RECT 70.415 58.4 70.635 59.16 ;
    RECT 71.115 58.4 71.335 59.16 ;
    RECT 71.815 58.4 72.035 59.16 ;
    RECT 72.515 58.4 72.735 59.16 ;
    RECT 73.215 58.4 73.435 59.16 ;
    RECT 73.915 58.4 74.835 59.16 ;
    RECT 75.315 58.4 75.535 59.16 ;
    RECT 76.015 58.4 76.225 59.16 ;
    RECT 76.705 58.4 76.92 59.16 ;
    RECT 77.4 58.4 77.62 59.16 ;
    RECT 78.1 58.4 78.32 59.16 ;
    RECT 78.8 58.4 79.02 59.16 ;
    RECT 79.5 58.4 81.115 59.16 ;
    RECT 81.595 58.4 81.815 59.16 ;
    RECT 82.295 58.4 82.515 59.16 ;
    RECT 82.995 58.4 83.055 59.16 ;
    RECT 83.055 58.31 83.335 59.25 ;
    RECT 83.335 58.4 83.505 59.16 ;
    RECT 26.71 57.64 26.88 58.4 ;
    RECT 26.88 57.55 27.16 58.49 ;
    RECT 27.16 57.64 27.32 58.4 ;
    RECT 27.8 57.64 28.02 58.4 ;
    RECT 28.5 57.64 28.72 58.4 ;
    RECT 29.2 57.64 30.815 58.4 ;
    RECT 31.295 57.64 31.515 58.4 ;
    RECT 31.995 57.64 32.21 58.4 ;
    RECT 32.69 57.64 32.91 58.4 ;
    RECT 33.39 57.64 33.61 58.4 ;
    RECT 34.09 57.64 34.31 58.4 ;
    RECT 34.79 57.64 35.005 58.4 ;
    RECT 35.485 57.64 36.405 58.4 ;
    RECT 36.885 57.64 37.105 58.4 ;
    RECT 37.585 57.64 37.8 58.4 ;
    RECT 38.28 57.64 38.5 58.4 ;
    RECT 38.98 57.64 39.2 58.4 ;
    RECT 39.68 57.64 39.895 58.4 ;
    RECT 40.375 57.64 40.595 58.4 ;
    RECT 41.075 57.64 41.995 58.4 ;
    RECT 42.475 57.64 42.69 58.4 ;
    RECT 43.17 57.64 43.39 58.4 ;
    RECT 43.87 57.64 44.09 58.4 ;
    RECT 44.57 57.64 44.79 58.4 ;
    RECT 45.27 57.64 45.485 58.4 ;
    RECT 45.965 57.64 46.185 58.4 ;
    RECT 46.665 57.64 47.58 58.4 ;
    RECT 48.06 57.64 48.28 58.4 ;
    RECT 48.76 57.64 48.98 58.4 ;
    RECT 49.46 57.64 49.68 58.4 ;
    RECT 50.16 57.64 50.375 58.4 ;
    RECT 50.855 57.64 51.775 58.4 ;
    RECT 52.255 57.64 53.17 58.4 ;
    RECT 53.65 57.64 53.87 58.4 ;
    RECT 54.35 57.64 54.57 58.4 ;
    RECT 55.05 57.64 55.265 58.4 ;
    RECT 55.745 57.64 55.965 58.4 ;
    RECT 56.445 57.64 56.665 58.4 ;
    RECT 57.145 57.64 58.06 58.4 ;
    RECT 58.54 57.64 59.46 58.4 ;
    RECT 59.94 57.64 60.16 58.4 ;
    RECT 60.64 57.64 60.855 58.4 ;
    RECT 61.335 57.64 61.555 58.4 ;
    RECT 62.035 57.64 62.25 58.4 ;
    RECT 62.73 57.64 63.65 58.4 ;
    RECT 64.13 57.64 64.345 58.4 ;
    RECT 64.825 57.64 65.045 58.4 ;
    RECT 65.525 57.64 65.745 58.4 ;
    RECT 66.225 57.64 66.445 58.4 ;
    RECT 66.925 57.64 67.14 58.4 ;
    RECT 67.62 57.64 67.84 58.4 ;
    RECT 68.32 57.64 69.235 58.4 ;
    RECT 69.715 57.64 69.935 58.4 ;
    RECT 70.415 57.64 70.635 58.4 ;
    RECT 71.115 57.64 71.335 58.4 ;
    RECT 71.815 57.64 72.035 58.4 ;
    RECT 72.515 57.64 72.735 58.4 ;
    RECT 73.215 57.64 73.435 58.4 ;
    RECT 73.915 57.64 74.835 58.4 ;
    RECT 75.315 57.64 75.535 58.4 ;
    RECT 76.015 57.64 76.225 58.4 ;
    RECT 76.705 57.64 76.92 58.4 ;
    RECT 77.4 57.64 77.62 58.4 ;
    RECT 78.1 57.64 78.32 58.4 ;
    RECT 78.8 57.64 79.02 58.4 ;
    RECT 79.5 57.64 81.115 58.4 ;
    RECT 81.595 57.64 81.815 58.4 ;
    RECT 82.295 57.64 82.515 58.4 ;
    RECT 82.995 57.64 83.055 58.4 ;
    RECT 83.055 57.55 83.335 58.49 ;
    RECT 83.335 57.64 83.505 58.4 ;
    RECT 26.71 56.88 26.88 57.64 ;
    RECT 26.88 56.79 27.16 57.73 ;
    RECT 27.16 56.88 27.32 57.64 ;
    RECT 27.8 56.88 28.02 57.64 ;
    RECT 28.5 56.88 28.72 57.64 ;
    RECT 29.2 56.88 30.815 57.64 ;
    RECT 31.295 56.88 31.515 57.64 ;
    RECT 31.995 56.88 32.21 57.64 ;
    RECT 32.69 56.88 32.91 57.64 ;
    RECT 33.39 56.88 33.61 57.64 ;
    RECT 34.09 56.88 34.31 57.64 ;
    RECT 34.79 56.88 35.005 57.64 ;
    RECT 35.485 56.88 36.405 57.64 ;
    RECT 36.885 56.88 37.105 57.64 ;
    RECT 37.585 56.88 37.8 57.64 ;
    RECT 38.28 56.88 38.5 57.64 ;
    RECT 38.98 56.88 39.2 57.64 ;
    RECT 39.68 56.88 39.895 57.64 ;
    RECT 40.375 56.88 40.595 57.64 ;
    RECT 41.075 56.88 41.995 57.64 ;
    RECT 42.475 56.88 42.69 57.64 ;
    RECT 43.17 56.88 43.39 57.64 ;
    RECT 43.87 56.88 44.09 57.64 ;
    RECT 44.57 56.88 44.79 57.64 ;
    RECT 45.27 56.88 45.485 57.64 ;
    RECT 45.965 56.88 46.185 57.64 ;
    RECT 46.665 56.88 47.58 57.64 ;
    RECT 48.06 56.88 48.28 57.64 ;
    RECT 48.76 56.88 48.98 57.64 ;
    RECT 49.46 56.88 49.68 57.64 ;
    RECT 50.16 56.88 50.375 57.64 ;
    RECT 50.855 56.88 51.775 57.64 ;
    RECT 52.255 56.88 53.17 57.64 ;
    RECT 53.65 56.88 53.87 57.64 ;
    RECT 54.35 56.88 54.57 57.64 ;
    RECT 55.05 56.88 55.265 57.64 ;
    RECT 55.745 56.88 55.965 57.64 ;
    RECT 56.445 56.88 56.665 57.64 ;
    RECT 57.145 56.88 58.06 57.64 ;
    RECT 58.54 56.88 59.46 57.64 ;
    RECT 59.94 56.88 60.16 57.64 ;
    RECT 60.64 56.88 60.855 57.64 ;
    RECT 61.335 56.88 61.555 57.64 ;
    RECT 62.035 56.88 62.25 57.64 ;
    RECT 62.73 56.88 63.65 57.64 ;
    RECT 64.13 56.88 64.345 57.64 ;
    RECT 64.825 56.88 65.045 57.64 ;
    RECT 65.525 56.88 65.745 57.64 ;
    RECT 66.225 56.88 66.445 57.64 ;
    RECT 66.925 56.88 67.14 57.64 ;
    RECT 67.62 56.88 67.84 57.64 ;
    RECT 68.32 56.88 69.235 57.64 ;
    RECT 69.715 56.88 69.935 57.64 ;
    RECT 70.415 56.88 70.635 57.64 ;
    RECT 71.115 56.88 71.335 57.64 ;
    RECT 71.815 56.88 72.035 57.64 ;
    RECT 72.515 56.88 72.735 57.64 ;
    RECT 73.215 56.88 73.435 57.64 ;
    RECT 73.915 56.88 74.835 57.64 ;
    RECT 75.315 56.88 75.535 57.64 ;
    RECT 76.015 56.88 76.225 57.64 ;
    RECT 76.705 56.88 76.92 57.64 ;
    RECT 77.4 56.88 77.62 57.64 ;
    RECT 78.1 56.88 78.32 57.64 ;
    RECT 78.8 56.88 79.02 57.64 ;
    RECT 79.5 56.88 81.115 57.64 ;
    RECT 81.595 56.88 81.815 57.64 ;
    RECT 82.295 56.88 82.515 57.64 ;
    RECT 82.995 56.88 83.055 57.64 ;
    RECT 83.055 56.79 83.335 57.73 ;
    RECT 83.335 56.88 83.505 57.64 ;
    RECT 26.71 56.12 26.88 56.88 ;
    RECT 26.88 56.03 27.16 56.97 ;
    RECT 27.16 56.12 27.32 56.88 ;
    RECT 27.8 56.12 28.02 56.88 ;
    RECT 28.5 56.12 28.72 56.88 ;
    RECT 29.2 56.12 30.815 56.88 ;
    RECT 31.295 56.12 31.515 56.88 ;
    RECT 31.995 56.12 32.21 56.88 ;
    RECT 32.69 56.12 32.91 56.88 ;
    RECT 33.39 56.12 33.61 56.88 ;
    RECT 34.09 56.12 34.31 56.88 ;
    RECT 34.79 56.12 35.005 56.88 ;
    RECT 35.485 56.12 36.405 56.88 ;
    RECT 36.885 56.12 37.105 56.88 ;
    RECT 37.585 56.12 37.8 56.88 ;
    RECT 38.28 56.12 38.5 56.88 ;
    RECT 38.98 56.12 39.2 56.88 ;
    RECT 39.68 56.12 39.895 56.88 ;
    RECT 40.375 56.12 40.595 56.88 ;
    RECT 41.075 56.12 41.995 56.88 ;
    RECT 42.475 56.12 42.69 56.88 ;
    RECT 43.17 56.12 43.39 56.88 ;
    RECT 43.87 56.12 44.09 56.88 ;
    RECT 44.57 56.12 44.79 56.88 ;
    RECT 45.27 56.12 45.485 56.88 ;
    RECT 45.965 56.12 46.185 56.88 ;
    RECT 46.665 56.12 47.58 56.88 ;
    RECT 48.06 56.12 48.28 56.88 ;
    RECT 48.76 56.12 48.98 56.88 ;
    RECT 49.46 56.12 49.68 56.88 ;
    RECT 50.16 56.12 50.375 56.88 ;
    RECT 50.855 56.12 51.775 56.88 ;
    RECT 52.255 56.12 53.17 56.88 ;
    RECT 53.65 56.12 53.87 56.88 ;
    RECT 54.35 56.12 54.57 56.88 ;
    RECT 55.05 56.12 55.265 56.88 ;
    RECT 55.745 56.12 55.965 56.88 ;
    RECT 56.445 56.12 56.665 56.88 ;
    RECT 57.145 56.12 58.06 56.88 ;
    RECT 58.54 56.12 59.46 56.88 ;
    RECT 59.94 56.12 60.16 56.88 ;
    RECT 60.64 56.12 60.855 56.88 ;
    RECT 61.335 56.12 61.555 56.88 ;
    RECT 62.035 56.12 62.25 56.88 ;
    RECT 62.73 56.12 63.65 56.88 ;
    RECT 64.13 56.12 64.345 56.88 ;
    RECT 64.825 56.12 65.045 56.88 ;
    RECT 65.525 56.12 65.745 56.88 ;
    RECT 66.225 56.12 66.445 56.88 ;
    RECT 66.925 56.12 67.14 56.88 ;
    RECT 67.62 56.12 67.84 56.88 ;
    RECT 68.32 56.12 69.235 56.88 ;
    RECT 69.715 56.12 69.935 56.88 ;
    RECT 70.415 56.12 70.635 56.88 ;
    RECT 71.115 56.12 71.335 56.88 ;
    RECT 71.815 56.12 72.035 56.88 ;
    RECT 72.515 56.12 72.735 56.88 ;
    RECT 73.215 56.12 73.435 56.88 ;
    RECT 73.915 56.12 74.835 56.88 ;
    RECT 75.315 56.12 75.535 56.88 ;
    RECT 76.015 56.12 76.225 56.88 ;
    RECT 76.705 56.12 76.92 56.88 ;
    RECT 77.4 56.12 77.62 56.88 ;
    RECT 78.1 56.12 78.32 56.88 ;
    RECT 78.8 56.12 79.02 56.88 ;
    RECT 79.5 56.12 81.115 56.88 ;
    RECT 81.595 56.12 81.815 56.88 ;
    RECT 82.295 56.12 82.515 56.88 ;
    RECT 82.995 56.12 83.055 56.88 ;
    RECT 83.055 56.03 83.335 56.97 ;
    RECT 83.335 56.12 83.505 56.88 ;
    RECT 26.71 55.36 26.88 56.12 ;
    RECT 26.88 55.27 27.16 56.21 ;
    RECT 27.16 55.36 27.32 56.12 ;
    RECT 27.8 55.36 28.02 56.12 ;
    RECT 28.5 55.36 28.72 56.12 ;
    RECT 29.2 55.36 30.815 56.12 ;
    RECT 31.295 55.36 31.515 56.12 ;
    RECT 31.995 55.36 32.21 56.12 ;
    RECT 32.69 55.36 32.91 56.12 ;
    RECT 33.39 55.36 33.61 56.12 ;
    RECT 34.09 55.36 34.31 56.12 ;
    RECT 34.79 55.36 35.005 56.12 ;
    RECT 35.485 55.36 36.405 56.12 ;
    RECT 36.885 55.36 37.105 56.12 ;
    RECT 37.585 55.36 37.8 56.12 ;
    RECT 38.28 55.36 38.5 56.12 ;
    RECT 38.98 55.36 39.2 56.12 ;
    RECT 39.68 55.36 39.895 56.12 ;
    RECT 40.375 55.36 40.595 56.12 ;
    RECT 41.075 55.36 41.995 56.12 ;
    RECT 42.475 55.36 42.69 56.12 ;
    RECT 43.17 55.36 43.39 56.12 ;
    RECT 43.87 55.36 44.09 56.12 ;
    RECT 44.57 55.36 44.79 56.12 ;
    RECT 45.27 55.36 45.485 56.12 ;
    RECT 45.965 55.36 46.185 56.12 ;
    RECT 46.665 55.36 47.58 56.12 ;
    RECT 48.06 55.36 48.28 56.12 ;
    RECT 48.76 55.36 48.98 56.12 ;
    RECT 49.46 55.36 49.68 56.12 ;
    RECT 50.16 55.36 50.375 56.12 ;
    RECT 50.855 55.36 51.775 56.12 ;
    RECT 52.255 55.36 53.17 56.12 ;
    RECT 53.65 55.36 53.87 56.12 ;
    RECT 54.35 55.36 54.57 56.12 ;
    RECT 55.05 55.36 55.265 56.12 ;
    RECT 55.745 55.36 55.965 56.12 ;
    RECT 56.445 55.36 56.665 56.12 ;
    RECT 57.145 55.36 58.06 56.12 ;
    RECT 58.54 55.36 59.46 56.12 ;
    RECT 59.94 55.36 60.16 56.12 ;
    RECT 60.64 55.36 60.855 56.12 ;
    RECT 61.335 55.36 61.555 56.12 ;
    RECT 62.035 55.36 62.25 56.12 ;
    RECT 62.73 55.36 63.65 56.12 ;
    RECT 64.13 55.36 64.345 56.12 ;
    RECT 64.825 55.36 65.045 56.12 ;
    RECT 65.525 55.36 65.745 56.12 ;
    RECT 66.225 55.36 66.445 56.12 ;
    RECT 66.925 55.36 67.14 56.12 ;
    RECT 67.62 55.36 67.84 56.12 ;
    RECT 68.32 55.36 69.235 56.12 ;
    RECT 69.715 55.36 69.935 56.12 ;
    RECT 70.415 55.36 70.635 56.12 ;
    RECT 71.115 55.36 71.335 56.12 ;
    RECT 71.815 55.36 72.035 56.12 ;
    RECT 72.515 55.36 72.735 56.12 ;
    RECT 73.215 55.36 73.435 56.12 ;
    RECT 73.915 55.36 74.835 56.12 ;
    RECT 75.315 55.36 75.535 56.12 ;
    RECT 76.015 55.36 76.225 56.12 ;
    RECT 76.705 55.36 76.92 56.12 ;
    RECT 77.4 55.36 77.62 56.12 ;
    RECT 78.1 55.36 78.32 56.12 ;
    RECT 78.8 55.36 79.02 56.12 ;
    RECT 79.5 55.36 81.115 56.12 ;
    RECT 81.595 55.36 81.815 56.12 ;
    RECT 82.295 55.36 82.515 56.12 ;
    RECT 82.995 55.36 83.055 56.12 ;
    RECT 83.055 55.27 83.335 56.21 ;
    RECT 83.335 55.36 83.505 56.12 ;
    RECT 26.71 54.6 26.88 55.36 ;
    RECT 26.88 54.51 27.16 55.45 ;
    RECT 27.16 54.6 27.32 55.36 ;
    RECT 27.8 54.6 28.02 55.36 ;
    RECT 28.5 54.6 28.72 55.36 ;
    RECT 29.2 54.6 30.815 55.36 ;
    RECT 31.295 54.6 31.515 55.36 ;
    RECT 31.995 54.6 32.21 55.36 ;
    RECT 32.69 54.6 32.91 55.36 ;
    RECT 33.39 54.6 33.61 55.36 ;
    RECT 34.09 54.6 34.31 55.36 ;
    RECT 34.79 54.6 35.005 55.36 ;
    RECT 35.485 54.6 36.405 55.36 ;
    RECT 36.885 54.6 37.105 55.36 ;
    RECT 37.585 54.6 37.8 55.36 ;
    RECT 38.28 54.6 38.5 55.36 ;
    RECT 38.98 54.6 39.2 55.36 ;
    RECT 39.68 54.6 39.895 55.36 ;
    RECT 40.375 54.6 40.595 55.36 ;
    RECT 41.075 54.6 41.995 55.36 ;
    RECT 42.475 54.6 42.69 55.36 ;
    RECT 43.17 54.6 43.39 55.36 ;
    RECT 43.87 54.6 44.09 55.36 ;
    RECT 44.57 54.6 44.79 55.36 ;
    RECT 45.27 54.6 45.485 55.36 ;
    RECT 45.965 54.6 46.185 55.36 ;
    RECT 46.665 54.6 47.58 55.36 ;
    RECT 48.06 54.6 48.28 55.36 ;
    RECT 48.76 54.6 48.98 55.36 ;
    RECT 49.46 54.6 49.68 55.36 ;
    RECT 50.16 54.6 50.375 55.36 ;
    RECT 50.855 54.6 51.775 55.36 ;
    RECT 52.255 54.6 53.17 55.36 ;
    RECT 53.65 54.6 53.87 55.36 ;
    RECT 54.35 54.6 54.57 55.36 ;
    RECT 55.05 54.6 55.265 55.36 ;
    RECT 55.745 54.6 55.965 55.36 ;
    RECT 56.445 54.6 56.665 55.36 ;
    RECT 57.145 54.6 58.06 55.36 ;
    RECT 58.54 54.6 59.46 55.36 ;
    RECT 59.94 54.6 60.16 55.36 ;
    RECT 60.64 54.6 60.855 55.36 ;
    RECT 61.335 54.6 61.555 55.36 ;
    RECT 62.035 54.6 62.25 55.36 ;
    RECT 62.73 54.6 63.65 55.36 ;
    RECT 64.13 54.6 64.345 55.36 ;
    RECT 64.825 54.6 65.045 55.36 ;
    RECT 65.525 54.6 65.745 55.36 ;
    RECT 66.225 54.6 66.445 55.36 ;
    RECT 66.925 54.6 67.14 55.36 ;
    RECT 67.62 54.6 67.84 55.36 ;
    RECT 68.32 54.6 69.235 55.36 ;
    RECT 69.715 54.6 69.935 55.36 ;
    RECT 70.415 54.6 70.635 55.36 ;
    RECT 71.115 54.6 71.335 55.36 ;
    RECT 71.815 54.6 72.035 55.36 ;
    RECT 72.515 54.6 72.735 55.36 ;
    RECT 73.215 54.6 73.435 55.36 ;
    RECT 73.915 54.6 74.835 55.36 ;
    RECT 75.315 54.6 75.535 55.36 ;
    RECT 76.015 54.6 76.225 55.36 ;
    RECT 76.705 54.6 76.92 55.36 ;
    RECT 77.4 54.6 77.62 55.36 ;
    RECT 78.1 54.6 78.32 55.36 ;
    RECT 78.8 54.6 79.02 55.36 ;
    RECT 79.5 54.6 81.115 55.36 ;
    RECT 81.595 54.6 81.815 55.36 ;
    RECT 82.295 54.6 82.515 55.36 ;
    RECT 82.995 54.6 83.055 55.36 ;
    RECT 83.055 54.51 83.335 55.45 ;
    RECT 83.335 54.6 83.505 55.36 ;
    RECT 26.71 53.84 26.88 54.6 ;
    RECT 26.88 53.75 27.16 54.69 ;
    RECT 27.16 53.84 27.32 54.6 ;
    RECT 27.8 53.84 28.02 54.6 ;
    RECT 28.5 53.84 28.72 54.6 ;
    RECT 29.2 53.84 30.815 54.6 ;
    RECT 31.295 53.84 31.515 54.6 ;
    RECT 31.995 53.84 32.21 54.6 ;
    RECT 32.69 53.84 32.91 54.6 ;
    RECT 33.39 53.84 33.61 54.6 ;
    RECT 34.09 53.84 34.31 54.6 ;
    RECT 34.79 53.84 35.005 54.6 ;
    RECT 35.485 53.84 36.405 54.6 ;
    RECT 36.885 53.84 37.105 54.6 ;
    RECT 37.585 53.84 37.8 54.6 ;
    RECT 38.28 53.84 38.5 54.6 ;
    RECT 38.98 53.84 39.2 54.6 ;
    RECT 39.68 53.84 39.895 54.6 ;
    RECT 40.375 53.84 40.595 54.6 ;
    RECT 41.075 53.84 41.995 54.6 ;
    RECT 42.475 53.84 42.69 54.6 ;
    RECT 43.17 53.84 43.39 54.6 ;
    RECT 43.87 53.84 44.09 54.6 ;
    RECT 44.57 53.84 44.79 54.6 ;
    RECT 45.27 53.84 45.485 54.6 ;
    RECT 45.965 53.84 46.185 54.6 ;
    RECT 46.665 53.84 47.58 54.6 ;
    RECT 48.06 53.84 48.28 54.6 ;
    RECT 48.76 53.84 48.98 54.6 ;
    RECT 49.46 53.84 49.68 54.6 ;
    RECT 50.16 53.84 50.375 54.6 ;
    RECT 50.855 53.84 51.775 54.6 ;
    RECT 52.255 53.84 53.17 54.6 ;
    RECT 53.65 53.84 53.87 54.6 ;
    RECT 54.35 53.84 54.57 54.6 ;
    RECT 55.05 53.84 55.265 54.6 ;
    RECT 55.745 53.84 55.965 54.6 ;
    RECT 56.445 53.84 56.665 54.6 ;
    RECT 57.145 53.84 58.06 54.6 ;
    RECT 58.54 53.84 59.46 54.6 ;
    RECT 59.94 53.84 60.16 54.6 ;
    RECT 60.64 53.84 60.855 54.6 ;
    RECT 61.335 53.84 61.555 54.6 ;
    RECT 62.035 53.84 62.25 54.6 ;
    RECT 62.73 53.84 63.65 54.6 ;
    RECT 64.13 53.84 64.345 54.6 ;
    RECT 64.825 53.84 65.045 54.6 ;
    RECT 65.525 53.84 65.745 54.6 ;
    RECT 66.225 53.84 66.445 54.6 ;
    RECT 66.925 53.84 67.14 54.6 ;
    RECT 67.62 53.84 67.84 54.6 ;
    RECT 68.32 53.84 69.235 54.6 ;
    RECT 69.715 53.84 69.935 54.6 ;
    RECT 70.415 53.84 70.635 54.6 ;
    RECT 71.115 53.84 71.335 54.6 ;
    RECT 71.815 53.84 72.035 54.6 ;
    RECT 72.515 53.84 72.735 54.6 ;
    RECT 73.215 53.84 73.435 54.6 ;
    RECT 73.915 53.84 74.835 54.6 ;
    RECT 75.315 53.84 75.535 54.6 ;
    RECT 76.015 53.84 76.225 54.6 ;
    RECT 76.705 53.84 76.92 54.6 ;
    RECT 77.4 53.84 77.62 54.6 ;
    RECT 78.1 53.84 78.32 54.6 ;
    RECT 78.8 53.84 79.02 54.6 ;
    RECT 79.5 53.84 81.115 54.6 ;
    RECT 81.595 53.84 81.815 54.6 ;
    RECT 82.295 53.84 82.515 54.6 ;
    RECT 82.995 53.84 83.055 54.6 ;
    RECT 83.055 53.75 83.335 54.69 ;
    RECT 83.335 53.84 83.505 54.6 ;
    RECT 26.71 53.08 26.88 53.84 ;
    RECT 26.88 52.99 27.16 53.93 ;
    RECT 27.16 53.08 27.32 53.84 ;
    RECT 27.8 53.08 28.02 53.84 ;
    RECT 28.5 53.08 28.72 53.84 ;
    RECT 29.2 53.08 30.815 53.84 ;
    RECT 31.295 53.08 31.515 53.84 ;
    RECT 31.995 53.08 32.21 53.84 ;
    RECT 32.69 53.08 32.91 53.84 ;
    RECT 33.39 53.08 33.61 53.84 ;
    RECT 34.09 53.08 34.31 53.84 ;
    RECT 34.79 53.08 35.005 53.84 ;
    RECT 35.485 53.08 36.405 53.84 ;
    RECT 36.885 53.08 37.105 53.84 ;
    RECT 37.585 53.08 37.8 53.84 ;
    RECT 38.28 53.08 38.5 53.84 ;
    RECT 38.98 53.08 39.2 53.84 ;
    RECT 39.68 53.08 39.895 53.84 ;
    RECT 40.375 53.08 40.595 53.84 ;
    RECT 41.075 53.08 41.995 53.84 ;
    RECT 42.475 53.08 42.69 53.84 ;
    RECT 43.17 53.08 43.39 53.84 ;
    RECT 43.87 53.08 44.09 53.84 ;
    RECT 44.57 53.08 44.79 53.84 ;
    RECT 45.27 53.08 45.485 53.84 ;
    RECT 45.965 53.08 46.185 53.84 ;
    RECT 46.665 53.08 47.58 53.84 ;
    RECT 48.06 53.08 48.28 53.84 ;
    RECT 48.76 53.08 48.98 53.84 ;
    RECT 49.46 53.08 49.68 53.84 ;
    RECT 50.16 53.08 50.375 53.84 ;
    RECT 50.855 53.08 51.775 53.84 ;
    RECT 52.255 53.08 53.17 53.84 ;
    RECT 53.65 53.08 53.87 53.84 ;
    RECT 54.35 53.08 54.57 53.84 ;
    RECT 55.05 53.08 55.265 53.84 ;
    RECT 55.745 53.08 55.965 53.84 ;
    RECT 56.445 53.08 56.665 53.84 ;
    RECT 57.145 53.08 58.06 53.84 ;
    RECT 58.54 53.08 59.46 53.84 ;
    RECT 59.94 53.08 60.16 53.84 ;
    RECT 60.64 53.08 60.855 53.84 ;
    RECT 61.335 53.08 61.555 53.84 ;
    RECT 62.035 53.08 62.25 53.84 ;
    RECT 62.73 53.08 63.65 53.84 ;
    RECT 64.13 53.08 64.345 53.84 ;
    RECT 64.825 53.08 65.045 53.84 ;
    RECT 65.525 53.08 65.745 53.84 ;
    RECT 66.225 53.08 66.445 53.84 ;
    RECT 66.925 53.08 67.14 53.84 ;
    RECT 67.62 53.08 67.84 53.84 ;
    RECT 68.32 53.08 69.235 53.84 ;
    RECT 69.715 53.08 69.935 53.84 ;
    RECT 70.415 53.08 70.635 53.84 ;
    RECT 71.115 53.08 71.335 53.84 ;
    RECT 71.815 53.08 72.035 53.84 ;
    RECT 72.515 53.08 72.735 53.84 ;
    RECT 73.215 53.08 73.435 53.84 ;
    RECT 73.915 53.08 74.835 53.84 ;
    RECT 75.315 53.08 75.535 53.84 ;
    RECT 76.015 53.08 76.225 53.84 ;
    RECT 76.705 53.08 76.92 53.84 ;
    RECT 77.4 53.08 77.62 53.84 ;
    RECT 78.1 53.08 78.32 53.84 ;
    RECT 78.8 53.08 79.02 53.84 ;
    RECT 79.5 53.08 81.115 53.84 ;
    RECT 81.595 53.08 81.815 53.84 ;
    RECT 82.295 53.08 82.515 53.84 ;
    RECT 82.995 53.08 83.055 53.84 ;
    RECT 83.055 52.99 83.335 53.93 ;
    RECT 83.335 53.08 83.505 53.84 ;
    RECT 26.71 52.32 26.88 53.08 ;
    RECT 26.88 52.23 27.16 53.17 ;
    RECT 27.16 52.32 27.32 53.08 ;
    RECT 27.8 52.32 28.02 53.08 ;
    RECT 28.5 52.32 28.72 53.08 ;
    RECT 29.2 52.32 30.815 53.08 ;
    RECT 31.295 52.32 31.515 53.08 ;
    RECT 31.995 52.32 32.21 53.08 ;
    RECT 32.69 52.32 32.91 53.08 ;
    RECT 33.39 52.32 33.61 53.08 ;
    RECT 34.09 52.32 34.31 53.08 ;
    RECT 34.79 52.32 35.005 53.08 ;
    RECT 35.485 52.32 36.405 53.08 ;
    RECT 36.885 52.32 37.105 53.08 ;
    RECT 37.585 52.32 37.8 53.08 ;
    RECT 38.28 52.32 38.5 53.08 ;
    RECT 38.98 52.32 39.2 53.08 ;
    RECT 39.68 52.32 39.895 53.08 ;
    RECT 40.375 52.32 40.595 53.08 ;
    RECT 41.075 52.32 41.995 53.08 ;
    RECT 42.475 52.32 42.69 53.08 ;
    RECT 43.17 52.32 43.39 53.08 ;
    RECT 43.87 52.32 44.09 53.08 ;
    RECT 44.57 52.32 44.79 53.08 ;
    RECT 45.27 52.32 45.485 53.08 ;
    RECT 45.965 52.32 46.185 53.08 ;
    RECT 46.665 52.32 47.58 53.08 ;
    RECT 48.06 52.32 48.28 53.08 ;
    RECT 48.76 52.32 48.98 53.08 ;
    RECT 49.46 52.32 49.68 53.08 ;
    RECT 50.16 52.32 50.375 53.08 ;
    RECT 50.855 52.32 51.775 53.08 ;
    RECT 52.255 52.32 53.17 53.08 ;
    RECT 53.65 52.32 53.87 53.08 ;
    RECT 54.35 52.32 54.57 53.08 ;
    RECT 55.05 52.32 55.265 53.08 ;
    RECT 55.745 52.32 55.965 53.08 ;
    RECT 56.445 52.32 56.665 53.08 ;
    RECT 57.145 52.32 58.06 53.08 ;
    RECT 58.54 52.32 59.46 53.08 ;
    RECT 59.94 52.32 60.16 53.08 ;
    RECT 60.64 52.32 60.855 53.08 ;
    RECT 61.335 52.32 61.555 53.08 ;
    RECT 62.035 52.32 62.25 53.08 ;
    RECT 62.73 52.32 63.65 53.08 ;
    RECT 64.13 52.32 64.345 53.08 ;
    RECT 64.825 52.32 65.045 53.08 ;
    RECT 65.525 52.32 65.745 53.08 ;
    RECT 66.225 52.32 66.445 53.08 ;
    RECT 66.925 52.32 67.14 53.08 ;
    RECT 67.62 52.32 67.84 53.08 ;
    RECT 68.32 52.32 69.235 53.08 ;
    RECT 69.715 52.32 69.935 53.08 ;
    RECT 70.415 52.32 70.635 53.08 ;
    RECT 71.115 52.32 71.335 53.08 ;
    RECT 71.815 52.32 72.035 53.08 ;
    RECT 72.515 52.32 72.735 53.08 ;
    RECT 73.215 52.32 73.435 53.08 ;
    RECT 73.915 52.32 74.835 53.08 ;
    RECT 75.315 52.32 75.535 53.08 ;
    RECT 76.015 52.32 76.225 53.08 ;
    RECT 76.705 52.32 76.92 53.08 ;
    RECT 77.4 52.32 77.62 53.08 ;
    RECT 78.1 52.32 78.32 53.08 ;
    RECT 78.8 52.32 79.02 53.08 ;
    RECT 79.5 52.32 81.115 53.08 ;
    RECT 81.595 52.32 81.815 53.08 ;
    RECT 82.295 52.32 82.515 53.08 ;
    RECT 82.995 52.32 83.055 53.08 ;
    RECT 83.055 52.23 83.335 53.17 ;
    RECT 83.335 52.32 83.505 53.08 ;
    RECT 26.71 51.56 26.88 52.32 ;
    RECT 26.88 51.47 27.16 52.41 ;
    RECT 27.16 51.56 27.32 52.32 ;
    RECT 27.8 51.56 28.02 52.32 ;
    RECT 28.5 51.56 28.72 52.32 ;
    RECT 29.2 51.56 30.815 52.32 ;
    RECT 31.295 51.56 31.515 52.32 ;
    RECT 31.995 51.56 32.21 52.32 ;
    RECT 32.69 51.56 32.91 52.32 ;
    RECT 33.39 51.56 33.61 52.32 ;
    RECT 34.09 51.56 34.31 52.32 ;
    RECT 34.79 51.56 35.005 52.32 ;
    RECT 35.485 51.56 36.405 52.32 ;
    RECT 36.885 51.56 37.105 52.32 ;
    RECT 37.585 51.56 37.8 52.32 ;
    RECT 38.28 51.56 38.5 52.32 ;
    RECT 38.98 51.56 39.2 52.32 ;
    RECT 39.68 51.56 39.895 52.32 ;
    RECT 40.375 51.56 40.595 52.32 ;
    RECT 41.075 51.56 41.995 52.32 ;
    RECT 42.475 51.56 42.69 52.32 ;
    RECT 43.17 51.56 43.39 52.32 ;
    RECT 43.87 51.56 44.09 52.32 ;
    RECT 44.57 51.56 44.79 52.32 ;
    RECT 45.27 51.56 45.485 52.32 ;
    RECT 45.965 51.56 46.185 52.32 ;
    RECT 46.665 51.56 47.58 52.32 ;
    RECT 48.06 51.56 48.28 52.32 ;
    RECT 48.76 51.56 48.98 52.32 ;
    RECT 49.46 51.56 49.68 52.32 ;
    RECT 50.16 51.56 50.375 52.32 ;
    RECT 50.855 51.56 51.775 52.32 ;
    RECT 52.255 51.56 53.17 52.32 ;
    RECT 53.65 51.56 53.87 52.32 ;
    RECT 54.35 51.56 54.57 52.32 ;
    RECT 55.05 51.56 55.265 52.32 ;
    RECT 55.745 51.56 55.965 52.32 ;
    RECT 56.445 51.56 56.665 52.32 ;
    RECT 57.145 51.56 58.06 52.32 ;
    RECT 58.54 51.56 59.46 52.32 ;
    RECT 59.94 51.56 60.16 52.32 ;
    RECT 60.64 51.56 60.855 52.32 ;
    RECT 61.335 51.56 61.555 52.32 ;
    RECT 62.035 51.56 62.25 52.32 ;
    RECT 62.73 51.56 63.65 52.32 ;
    RECT 64.13 51.56 64.345 52.32 ;
    RECT 64.825 51.56 65.045 52.32 ;
    RECT 65.525 51.56 65.745 52.32 ;
    RECT 66.225 51.56 66.445 52.32 ;
    RECT 66.925 51.56 67.14 52.32 ;
    RECT 67.62 51.56 67.84 52.32 ;
    RECT 68.32 51.56 69.235 52.32 ;
    RECT 69.715 51.56 69.935 52.32 ;
    RECT 70.415 51.56 70.635 52.32 ;
    RECT 71.115 51.56 71.335 52.32 ;
    RECT 71.815 51.56 72.035 52.32 ;
    RECT 72.515 51.56 72.735 52.32 ;
    RECT 73.215 51.56 73.435 52.32 ;
    RECT 73.915 51.56 74.835 52.32 ;
    RECT 75.315 51.56 75.535 52.32 ;
    RECT 76.015 51.56 76.225 52.32 ;
    RECT 76.705 51.56 76.92 52.32 ;
    RECT 77.4 51.56 77.62 52.32 ;
    RECT 78.1 51.56 78.32 52.32 ;
    RECT 78.8 51.56 79.02 52.32 ;
    RECT 79.5 51.56 81.115 52.32 ;
    RECT 81.595 51.56 81.815 52.32 ;
    RECT 82.295 51.56 82.515 52.32 ;
    RECT 82.995 51.56 83.055 52.32 ;
    RECT 83.055 51.47 83.335 52.41 ;
    RECT 83.335 51.56 83.505 52.32 ;
    RECT 26.71 50.8 26.88 51.56 ;
    RECT 26.88 50.71 27.16 51.65 ;
    RECT 27.16 50.8 27.32 51.56 ;
    RECT 27.8 50.8 28.02 51.56 ;
    RECT 28.5 50.8 28.72 51.56 ;
    RECT 29.2 50.8 30.815 51.56 ;
    RECT 31.295 50.8 31.515 51.56 ;
    RECT 31.995 50.8 32.21 51.56 ;
    RECT 32.69 50.8 32.91 51.56 ;
    RECT 33.39 50.8 33.61 51.56 ;
    RECT 34.09 50.8 34.31 51.56 ;
    RECT 34.79 50.8 35.005 51.56 ;
    RECT 35.485 50.8 36.405 51.56 ;
    RECT 36.885 50.8 37.105 51.56 ;
    RECT 37.585 50.8 37.8 51.56 ;
    RECT 38.28 50.8 38.5 51.56 ;
    RECT 38.98 50.8 39.2 51.56 ;
    RECT 39.68 50.8 39.895 51.56 ;
    RECT 40.375 50.8 40.595 51.56 ;
    RECT 41.075 50.8 41.995 51.56 ;
    RECT 42.475 50.8 42.69 51.56 ;
    RECT 43.17 50.8 43.39 51.56 ;
    RECT 43.87 50.8 44.09 51.56 ;
    RECT 44.57 50.8 44.79 51.56 ;
    RECT 45.27 50.8 45.485 51.56 ;
    RECT 45.965 50.8 46.185 51.56 ;
    RECT 46.665 50.8 47.58 51.56 ;
    RECT 48.06 50.8 48.28 51.56 ;
    RECT 48.76 50.8 48.98 51.56 ;
    RECT 49.46 50.8 49.68 51.56 ;
    RECT 50.16 50.8 50.375 51.56 ;
    RECT 50.855 50.8 51.775 51.56 ;
    RECT 52.255 50.8 53.17 51.56 ;
    RECT 53.65 50.8 53.87 51.56 ;
    RECT 54.35 50.8 54.57 51.56 ;
    RECT 55.05 50.8 55.265 51.56 ;
    RECT 55.745 50.8 55.965 51.56 ;
    RECT 56.445 50.8 56.665 51.56 ;
    RECT 57.145 50.8 58.06 51.56 ;
    RECT 58.54 50.8 59.46 51.56 ;
    RECT 59.94 50.8 60.16 51.56 ;
    RECT 60.64 50.8 60.855 51.56 ;
    RECT 61.335 50.8 61.555 51.56 ;
    RECT 62.035 50.8 62.25 51.56 ;
    RECT 62.73 50.8 63.65 51.56 ;
    RECT 64.13 50.8 64.345 51.56 ;
    RECT 64.825 50.8 65.045 51.56 ;
    RECT 65.525 50.8 65.745 51.56 ;
    RECT 66.225 50.8 66.445 51.56 ;
    RECT 66.925 50.8 67.14 51.56 ;
    RECT 67.62 50.8 67.84 51.56 ;
    RECT 68.32 50.8 69.235 51.56 ;
    RECT 69.715 50.8 69.935 51.56 ;
    RECT 70.415 50.8 70.635 51.56 ;
    RECT 71.115 50.8 71.335 51.56 ;
    RECT 71.815 50.8 72.035 51.56 ;
    RECT 72.515 50.8 72.735 51.56 ;
    RECT 73.215 50.8 73.435 51.56 ;
    RECT 73.915 50.8 74.835 51.56 ;
    RECT 75.315 50.8 75.535 51.56 ;
    RECT 76.015 50.8 76.225 51.56 ;
    RECT 76.705 50.8 76.92 51.56 ;
    RECT 77.4 50.8 77.62 51.56 ;
    RECT 78.1 50.8 78.32 51.56 ;
    RECT 78.8 50.8 79.02 51.56 ;
    RECT 79.5 50.8 81.115 51.56 ;
    RECT 81.595 50.8 81.815 51.56 ;
    RECT 82.295 50.8 82.515 51.56 ;
    RECT 82.995 50.8 83.055 51.56 ;
    RECT 83.055 50.71 83.335 51.65 ;
    RECT 83.335 50.8 83.505 51.56 ;
    RECT 26.71 50.04 26.88 50.8 ;
    RECT 26.88 49.95 27.16 50.89 ;
    RECT 27.16 50.04 27.32 50.8 ;
    RECT 27.8 50.04 28.02 50.8 ;
    RECT 28.5 50.04 28.72 50.8 ;
    RECT 29.2 50.04 30.815 50.8 ;
    RECT 31.295 50.04 31.515 50.8 ;
    RECT 31.995 50.04 32.21 50.8 ;
    RECT 32.69 50.04 32.91 50.8 ;
    RECT 33.39 50.04 33.61 50.8 ;
    RECT 34.09 50.04 34.31 50.8 ;
    RECT 34.79 50.04 35.005 50.8 ;
    RECT 35.485 50.04 36.405 50.8 ;
    RECT 36.885 50.04 37.105 50.8 ;
    RECT 37.585 50.04 37.8 50.8 ;
    RECT 38.28 50.04 38.5 50.8 ;
    RECT 38.98 50.04 39.2 50.8 ;
    RECT 39.68 50.04 39.895 50.8 ;
    RECT 40.375 50.04 40.595 50.8 ;
    RECT 41.075 50.04 41.995 50.8 ;
    RECT 42.475 50.04 42.69 50.8 ;
    RECT 43.17 50.04 43.39 50.8 ;
    RECT 43.87 50.04 44.09 50.8 ;
    RECT 44.57 50.04 44.79 50.8 ;
    RECT 45.27 50.04 45.485 50.8 ;
    RECT 45.965 50.04 46.185 50.8 ;
    RECT 46.665 50.04 47.58 50.8 ;
    RECT 48.06 50.04 48.28 50.8 ;
    RECT 48.76 50.04 48.98 50.8 ;
    RECT 49.46 50.04 49.68 50.8 ;
    RECT 50.16 50.04 50.375 50.8 ;
    RECT 50.855 50.04 51.775 50.8 ;
    RECT 52.255 50.04 53.17 50.8 ;
    RECT 53.65 50.04 53.87 50.8 ;
    RECT 54.35 50.04 54.57 50.8 ;
    RECT 55.05 50.04 55.265 50.8 ;
    RECT 55.745 50.04 55.965 50.8 ;
    RECT 56.445 50.04 56.665 50.8 ;
    RECT 57.145 50.04 58.06 50.8 ;
    RECT 58.54 50.04 59.46 50.8 ;
    RECT 59.94 50.04 60.16 50.8 ;
    RECT 60.64 50.04 60.855 50.8 ;
    RECT 61.335 50.04 61.555 50.8 ;
    RECT 62.035 50.04 62.25 50.8 ;
    RECT 62.73 50.04 63.65 50.8 ;
    RECT 64.13 50.04 64.345 50.8 ;
    RECT 64.825 50.04 65.045 50.8 ;
    RECT 65.525 50.04 65.745 50.8 ;
    RECT 66.225 50.04 66.445 50.8 ;
    RECT 66.925 50.04 67.14 50.8 ;
    RECT 67.62 50.04 67.84 50.8 ;
    RECT 68.32 50.04 69.235 50.8 ;
    RECT 69.715 50.04 69.935 50.8 ;
    RECT 70.415 50.04 70.635 50.8 ;
    RECT 71.115 50.04 71.335 50.8 ;
    RECT 71.815 50.04 72.035 50.8 ;
    RECT 72.515 50.04 72.735 50.8 ;
    RECT 73.215 50.04 73.435 50.8 ;
    RECT 73.915 50.04 74.835 50.8 ;
    RECT 75.315 50.04 75.535 50.8 ;
    RECT 76.015 50.04 76.225 50.8 ;
    RECT 76.705 50.04 76.92 50.8 ;
    RECT 77.4 50.04 77.62 50.8 ;
    RECT 78.1 50.04 78.32 50.8 ;
    RECT 78.8 50.04 79.02 50.8 ;
    RECT 79.5 50.04 81.115 50.8 ;
    RECT 81.595 50.04 81.815 50.8 ;
    RECT 82.295 50.04 82.515 50.8 ;
    RECT 82.995 50.04 83.055 50.8 ;
    RECT 83.055 49.95 83.335 50.89 ;
    RECT 83.335 50.04 83.505 50.8 ;
    RECT 26.71 49.28 26.88 50.04 ;
    RECT 26.88 49.19 27.16 50.13 ;
    RECT 27.16 49.28 27.32 50.04 ;
    RECT 27.8 49.28 28.02 50.04 ;
    RECT 28.5 49.28 28.72 50.04 ;
    RECT 29.2 49.28 30.815 50.04 ;
    RECT 31.295 49.28 31.515 50.04 ;
    RECT 31.995 49.28 32.21 50.04 ;
    RECT 32.69 49.28 32.91 50.04 ;
    RECT 33.39 49.28 33.61 50.04 ;
    RECT 34.09 49.28 34.31 50.04 ;
    RECT 34.79 49.28 35.005 50.04 ;
    RECT 35.485 49.28 36.405 50.04 ;
    RECT 36.885 49.28 37.105 50.04 ;
    RECT 37.585 49.28 37.8 50.04 ;
    RECT 38.28 49.28 38.5 50.04 ;
    RECT 38.98 49.28 39.2 50.04 ;
    RECT 39.68 49.28 39.895 50.04 ;
    RECT 40.375 49.28 40.595 50.04 ;
    RECT 41.075 49.28 41.995 50.04 ;
    RECT 42.475 49.28 42.69 50.04 ;
    RECT 43.17 49.28 43.39 50.04 ;
    RECT 43.87 49.28 44.09 50.04 ;
    RECT 44.57 49.28 44.79 50.04 ;
    RECT 45.27 49.28 45.485 50.04 ;
    RECT 45.965 49.28 46.185 50.04 ;
    RECT 46.665 49.28 47.58 50.04 ;
    RECT 48.06 49.28 48.28 50.04 ;
    RECT 48.76 49.28 48.98 50.04 ;
    RECT 49.46 49.28 49.68 50.04 ;
    RECT 50.16 49.28 50.375 50.04 ;
    RECT 50.855 49.28 51.775 50.04 ;
    RECT 52.255 49.28 53.17 50.04 ;
    RECT 53.65 49.28 53.87 50.04 ;
    RECT 54.35 49.28 54.57 50.04 ;
    RECT 55.05 49.28 55.265 50.04 ;
    RECT 55.745 49.28 55.965 50.04 ;
    RECT 56.445 49.28 56.665 50.04 ;
    RECT 57.145 49.28 58.06 50.04 ;
    RECT 58.54 49.28 59.46 50.04 ;
    RECT 59.94 49.28 60.16 50.04 ;
    RECT 60.64 49.28 60.855 50.04 ;
    RECT 61.335 49.28 61.555 50.04 ;
    RECT 62.035 49.28 62.25 50.04 ;
    RECT 62.73 49.28 63.65 50.04 ;
    RECT 64.13 49.28 64.345 50.04 ;
    RECT 64.825 49.28 65.045 50.04 ;
    RECT 65.525 49.28 65.745 50.04 ;
    RECT 66.225 49.28 66.445 50.04 ;
    RECT 66.925 49.28 67.14 50.04 ;
    RECT 67.62 49.28 67.84 50.04 ;
    RECT 68.32 49.28 69.235 50.04 ;
    RECT 69.715 49.28 69.935 50.04 ;
    RECT 70.415 49.28 70.635 50.04 ;
    RECT 71.115 49.28 71.335 50.04 ;
    RECT 71.815 49.28 72.035 50.04 ;
    RECT 72.515 49.28 72.735 50.04 ;
    RECT 73.215 49.28 73.435 50.04 ;
    RECT 73.915 49.28 74.835 50.04 ;
    RECT 75.315 49.28 75.535 50.04 ;
    RECT 76.015 49.28 76.225 50.04 ;
    RECT 76.705 49.28 76.92 50.04 ;
    RECT 77.4 49.28 77.62 50.04 ;
    RECT 78.1 49.28 78.32 50.04 ;
    RECT 78.8 49.28 79.02 50.04 ;
    RECT 79.5 49.28 81.115 50.04 ;
    RECT 81.595 49.28 81.815 50.04 ;
    RECT 82.295 49.28 82.515 50.04 ;
    RECT 82.995 49.28 83.055 50.04 ;
    RECT 83.055 49.19 83.335 50.13 ;
    RECT 83.335 49.28 83.505 50.04 ;
    RECT 26.71 48.52 26.88 49.28 ;
    RECT 26.88 48.43 27.16 49.37 ;
    RECT 27.16 48.52 27.32 49.28 ;
    RECT 27.8 48.52 28.02 49.28 ;
    RECT 28.5 48.52 28.72 49.28 ;
    RECT 29.2 48.52 30.815 49.28 ;
    RECT 31.295 48.52 31.515 49.28 ;
    RECT 31.995 48.52 32.21 49.28 ;
    RECT 32.69 48.52 32.91 49.28 ;
    RECT 33.39 48.52 33.61 49.28 ;
    RECT 34.09 48.52 34.31 49.28 ;
    RECT 34.79 48.52 35.005 49.28 ;
    RECT 35.485 48.52 36.405 49.28 ;
    RECT 36.885 48.52 37.105 49.28 ;
    RECT 37.585 48.52 37.8 49.28 ;
    RECT 38.28 48.52 38.5 49.28 ;
    RECT 38.98 48.52 39.2 49.28 ;
    RECT 39.68 48.52 39.895 49.28 ;
    RECT 40.375 48.52 40.595 49.28 ;
    RECT 41.075 48.52 41.995 49.28 ;
    RECT 42.475 48.52 42.69 49.28 ;
    RECT 43.17 48.52 43.39 49.28 ;
    RECT 43.87 48.52 44.09 49.28 ;
    RECT 44.57 48.52 44.79 49.28 ;
    RECT 45.27 48.52 45.485 49.28 ;
    RECT 45.965 48.52 46.185 49.28 ;
    RECT 46.665 48.52 47.58 49.28 ;
    RECT 48.06 48.52 48.28 49.28 ;
    RECT 48.76 48.52 48.98 49.28 ;
    RECT 49.46 48.52 49.68 49.28 ;
    RECT 50.16 48.52 50.375 49.28 ;
    RECT 50.855 48.52 51.775 49.28 ;
    RECT 52.255 48.52 53.17 49.28 ;
    RECT 53.65 48.52 53.87 49.28 ;
    RECT 54.35 48.52 54.57 49.28 ;
    RECT 55.05 48.52 55.265 49.28 ;
    RECT 55.745 48.52 55.965 49.28 ;
    RECT 56.445 48.52 56.665 49.28 ;
    RECT 57.145 48.52 58.06 49.28 ;
    RECT 58.54 48.52 59.46 49.28 ;
    RECT 59.94 48.52 60.16 49.28 ;
    RECT 60.64 48.52 60.855 49.28 ;
    RECT 61.335 48.52 61.555 49.28 ;
    RECT 62.035 48.52 62.25 49.28 ;
    RECT 62.73 48.52 63.65 49.28 ;
    RECT 64.13 48.52 64.345 49.28 ;
    RECT 64.825 48.52 65.045 49.28 ;
    RECT 65.525 48.52 65.745 49.28 ;
    RECT 66.225 48.52 66.445 49.28 ;
    RECT 66.925 48.52 67.14 49.28 ;
    RECT 67.62 48.52 67.84 49.28 ;
    RECT 68.32 48.52 69.235 49.28 ;
    RECT 69.715 48.52 69.935 49.28 ;
    RECT 70.415 48.52 70.635 49.28 ;
    RECT 71.115 48.52 71.335 49.28 ;
    RECT 71.815 48.52 72.035 49.28 ;
    RECT 72.515 48.52 72.735 49.28 ;
    RECT 73.215 48.52 73.435 49.28 ;
    RECT 73.915 48.52 74.835 49.28 ;
    RECT 75.315 48.52 75.535 49.28 ;
    RECT 76.015 48.52 76.225 49.28 ;
    RECT 76.705 48.52 76.92 49.28 ;
    RECT 77.4 48.52 77.62 49.28 ;
    RECT 78.1 48.52 78.32 49.28 ;
    RECT 78.8 48.52 79.02 49.28 ;
    RECT 79.5 48.52 81.115 49.28 ;
    RECT 81.595 48.52 81.815 49.28 ;
    RECT 82.295 48.52 82.515 49.28 ;
    RECT 82.995 48.52 83.055 49.28 ;
    RECT 83.055 48.43 83.335 49.37 ;
    RECT 83.335 48.52 83.505 49.28 ;
    RECT 26.71 47.76 26.88 48.52 ;
    RECT 26.88 47.67 27.16 48.61 ;
    RECT 27.16 47.76 27.32 48.52 ;
    RECT 27.8 47.76 28.02 48.52 ;
    RECT 28.5 47.76 28.72 48.52 ;
    RECT 29.2 47.76 30.815 48.52 ;
    RECT 31.295 47.76 31.515 48.52 ;
    RECT 31.995 47.76 32.21 48.52 ;
    RECT 32.69 47.76 32.91 48.52 ;
    RECT 33.39 47.76 33.61 48.52 ;
    RECT 34.09 47.76 34.31 48.52 ;
    RECT 34.79 47.76 35.005 48.52 ;
    RECT 35.485 47.76 36.405 48.52 ;
    RECT 36.885 47.76 37.105 48.52 ;
    RECT 37.585 47.76 37.8 48.52 ;
    RECT 38.28 47.76 38.5 48.52 ;
    RECT 38.98 47.76 39.2 48.52 ;
    RECT 39.68 47.76 39.895 48.52 ;
    RECT 40.375 47.76 40.595 48.52 ;
    RECT 41.075 47.76 41.995 48.52 ;
    RECT 42.475 47.76 42.69 48.52 ;
    RECT 43.17 47.76 43.39 48.52 ;
    RECT 43.87 47.76 44.09 48.52 ;
    RECT 44.57 47.76 44.79 48.52 ;
    RECT 45.27 47.76 45.485 48.52 ;
    RECT 45.965 47.76 46.185 48.52 ;
    RECT 46.665 47.76 47.58 48.52 ;
    RECT 48.06 47.76 48.28 48.52 ;
    RECT 48.76 47.76 48.98 48.52 ;
    RECT 49.46 47.76 49.68 48.52 ;
    RECT 50.16 47.76 50.375 48.52 ;
    RECT 50.855 47.76 51.775 48.52 ;
    RECT 52.255 47.76 53.17 48.52 ;
    RECT 53.65 47.76 53.87 48.52 ;
    RECT 54.35 47.76 54.57 48.52 ;
    RECT 55.05 47.76 55.265 48.52 ;
    RECT 55.745 47.76 55.965 48.52 ;
    RECT 56.445 47.76 56.665 48.52 ;
    RECT 57.145 47.76 58.06 48.52 ;
    RECT 58.54 47.76 59.46 48.52 ;
    RECT 59.94 47.76 60.16 48.52 ;
    RECT 60.64 47.76 60.855 48.52 ;
    RECT 61.335 47.76 61.555 48.52 ;
    RECT 62.035 47.76 62.25 48.52 ;
    RECT 62.73 47.76 63.65 48.52 ;
    RECT 64.13 47.76 64.345 48.52 ;
    RECT 64.825 47.76 65.045 48.52 ;
    RECT 65.525 47.76 65.745 48.52 ;
    RECT 66.225 47.76 66.445 48.52 ;
    RECT 66.925 47.76 67.14 48.52 ;
    RECT 67.62 47.76 67.84 48.52 ;
    RECT 68.32 47.76 69.235 48.52 ;
    RECT 69.715 47.76 69.935 48.52 ;
    RECT 70.415 47.76 70.635 48.52 ;
    RECT 71.115 47.76 71.335 48.52 ;
    RECT 71.815 47.76 72.035 48.52 ;
    RECT 72.515 47.76 72.735 48.52 ;
    RECT 73.215 47.76 73.435 48.52 ;
    RECT 73.915 47.76 74.835 48.52 ;
    RECT 75.315 47.76 75.535 48.52 ;
    RECT 76.015 47.76 76.225 48.52 ;
    RECT 76.705 47.76 76.92 48.52 ;
    RECT 77.4 47.76 77.62 48.52 ;
    RECT 78.1 47.76 78.32 48.52 ;
    RECT 78.8 47.76 79.02 48.52 ;
    RECT 79.5 47.76 81.115 48.52 ;
    RECT 81.595 47.76 81.815 48.52 ;
    RECT 82.295 47.76 82.515 48.52 ;
    RECT 82.995 47.76 83.055 48.52 ;
    RECT 83.055 47.67 83.335 48.61 ;
    RECT 83.335 47.76 83.505 48.52 ;
    RECT 26.71 47.0 26.88 47.76 ;
    RECT 26.88 46.91 27.16 47.85 ;
    RECT 27.16 47.0 27.32 47.76 ;
    RECT 27.8 47.0 28.02 47.76 ;
    RECT 28.5 47.0 28.72 47.76 ;
    RECT 29.2 47.0 30.815 47.76 ;
    RECT 31.295 47.0 31.515 47.76 ;
    RECT 31.995 47.0 32.21 47.76 ;
    RECT 32.69 47.0 32.91 47.76 ;
    RECT 33.39 47.0 33.61 47.76 ;
    RECT 34.09 47.0 34.31 47.76 ;
    RECT 34.79 47.0 35.005 47.76 ;
    RECT 35.485 47.0 36.405 47.76 ;
    RECT 36.885 47.0 37.105 47.76 ;
    RECT 37.585 47.0 37.8 47.76 ;
    RECT 38.28 47.0 38.5 47.76 ;
    RECT 38.98 47.0 39.2 47.76 ;
    RECT 39.68 47.0 39.895 47.76 ;
    RECT 40.375 47.0 40.595 47.76 ;
    RECT 41.075 47.0 41.995 47.76 ;
    RECT 42.475 47.0 42.69 47.76 ;
    RECT 43.17 47.0 43.39 47.76 ;
    RECT 43.87 47.0 44.09 47.76 ;
    RECT 44.57 47.0 44.79 47.76 ;
    RECT 45.27 47.0 45.485 47.76 ;
    RECT 45.965 47.0 46.185 47.76 ;
    RECT 46.665 47.0 47.58 47.76 ;
    RECT 48.06 47.0 48.28 47.76 ;
    RECT 48.76 47.0 48.98 47.76 ;
    RECT 49.46 47.0 49.68 47.76 ;
    RECT 50.16 47.0 50.375 47.76 ;
    RECT 50.855 47.0 51.775 47.76 ;
    RECT 52.255 47.0 53.17 47.76 ;
    RECT 53.65 47.0 53.87 47.76 ;
    RECT 54.35 47.0 54.57 47.76 ;
    RECT 55.05 47.0 55.265 47.76 ;
    RECT 55.745 47.0 55.965 47.76 ;
    RECT 56.445 47.0 56.665 47.76 ;
    RECT 57.145 47.0 58.06 47.76 ;
    RECT 58.54 47.0 59.46 47.76 ;
    RECT 59.94 47.0 60.16 47.76 ;
    RECT 60.64 47.0 60.855 47.76 ;
    RECT 61.335 47.0 61.555 47.76 ;
    RECT 62.035 47.0 62.25 47.76 ;
    RECT 62.73 47.0 63.65 47.76 ;
    RECT 64.13 47.0 64.345 47.76 ;
    RECT 64.825 47.0 65.045 47.76 ;
    RECT 65.525 47.0 65.745 47.76 ;
    RECT 66.225 47.0 66.445 47.76 ;
    RECT 66.925 47.0 67.14 47.76 ;
    RECT 67.62 47.0 67.84 47.76 ;
    RECT 68.32 47.0 69.235 47.76 ;
    RECT 69.715 47.0 69.935 47.76 ;
    RECT 70.415 47.0 70.635 47.76 ;
    RECT 71.115 47.0 71.335 47.76 ;
    RECT 71.815 47.0 72.035 47.76 ;
    RECT 72.515 47.0 72.735 47.76 ;
    RECT 73.215 47.0 73.435 47.76 ;
    RECT 73.915 47.0 74.835 47.76 ;
    RECT 75.315 47.0 75.535 47.76 ;
    RECT 76.015 47.0 76.225 47.76 ;
    RECT 76.705 47.0 76.92 47.76 ;
    RECT 77.4 47.0 77.62 47.76 ;
    RECT 78.1 47.0 78.32 47.76 ;
    RECT 78.8 47.0 79.02 47.76 ;
    RECT 79.5 47.0 81.115 47.76 ;
    RECT 81.595 47.0 81.815 47.76 ;
    RECT 82.295 47.0 82.515 47.76 ;
    RECT 82.995 47.0 83.055 47.76 ;
    RECT 83.055 46.91 83.335 47.85 ;
    RECT 83.335 47.0 83.505 47.76 ;
    RECT 26.71 46.24 26.88 47.0 ;
    RECT 26.88 46.15 27.16 47.09 ;
    RECT 27.16 46.24 27.32 47.0 ;
    RECT 27.8 46.24 28.02 47.0 ;
    RECT 28.5 46.24 28.72 47.0 ;
    RECT 29.2 46.24 30.815 47.0 ;
    RECT 31.295 46.24 31.515 47.0 ;
    RECT 31.995 46.24 32.21 47.0 ;
    RECT 32.69 46.24 32.91 47.0 ;
    RECT 33.39 46.24 33.61 47.0 ;
    RECT 34.09 46.24 34.31 47.0 ;
    RECT 34.79 46.24 35.005 47.0 ;
    RECT 35.485 46.24 36.405 47.0 ;
    RECT 36.885 46.24 37.105 47.0 ;
    RECT 37.585 46.24 37.8 47.0 ;
    RECT 38.28 46.24 38.5 47.0 ;
    RECT 38.98 46.24 39.2 47.0 ;
    RECT 39.68 46.24 39.895 47.0 ;
    RECT 40.375 46.24 40.595 47.0 ;
    RECT 41.075 46.24 41.995 47.0 ;
    RECT 42.475 46.24 42.69 47.0 ;
    RECT 43.17 46.24 43.39 47.0 ;
    RECT 43.87 46.24 44.09 47.0 ;
    RECT 44.57 46.24 44.79 47.0 ;
    RECT 45.27 46.24 45.485 47.0 ;
    RECT 45.965 46.24 46.185 47.0 ;
    RECT 46.665 46.24 47.58 47.0 ;
    RECT 48.06 46.24 48.28 47.0 ;
    RECT 48.76 46.24 48.98 47.0 ;
    RECT 49.46 46.24 49.68 47.0 ;
    RECT 50.16 46.24 50.375 47.0 ;
    RECT 50.855 46.24 51.775 47.0 ;
    RECT 52.255 46.24 53.17 47.0 ;
    RECT 53.65 46.24 53.87 47.0 ;
    RECT 54.35 46.24 54.57 47.0 ;
    RECT 55.05 46.24 55.265 47.0 ;
    RECT 55.745 46.24 55.965 47.0 ;
    RECT 56.445 46.24 56.665 47.0 ;
    RECT 57.145 46.24 58.06 47.0 ;
    RECT 58.54 46.24 59.46 47.0 ;
    RECT 59.94 46.24 60.16 47.0 ;
    RECT 60.64 46.24 60.855 47.0 ;
    RECT 61.335 46.24 61.555 47.0 ;
    RECT 62.035 46.24 62.25 47.0 ;
    RECT 62.73 46.24 63.65 47.0 ;
    RECT 64.13 46.24 64.345 47.0 ;
    RECT 64.825 46.24 65.045 47.0 ;
    RECT 65.525 46.24 65.745 47.0 ;
    RECT 66.225 46.24 66.445 47.0 ;
    RECT 66.925 46.24 67.14 47.0 ;
    RECT 67.62 46.24 67.84 47.0 ;
    RECT 68.32 46.24 69.235 47.0 ;
    RECT 69.715 46.24 69.935 47.0 ;
    RECT 70.415 46.24 70.635 47.0 ;
    RECT 71.115 46.24 71.335 47.0 ;
    RECT 71.815 46.24 72.035 47.0 ;
    RECT 72.515 46.24 72.735 47.0 ;
    RECT 73.215 46.24 73.435 47.0 ;
    RECT 73.915 46.24 74.835 47.0 ;
    RECT 75.315 46.24 75.535 47.0 ;
    RECT 76.015 46.24 76.225 47.0 ;
    RECT 76.705 46.24 76.92 47.0 ;
    RECT 77.4 46.24 77.62 47.0 ;
    RECT 78.1 46.24 78.32 47.0 ;
    RECT 78.8 46.24 79.02 47.0 ;
    RECT 79.5 46.24 81.115 47.0 ;
    RECT 81.595 46.24 81.815 47.0 ;
    RECT 82.295 46.24 82.515 47.0 ;
    RECT 82.995 46.24 83.055 47.0 ;
    RECT 83.055 46.15 83.335 47.09 ;
    RECT 83.335 46.24 83.505 47.0 ;
    RECT 26.71 45.48 26.88 46.24 ;
    RECT 26.88 45.39 27.16 46.33 ;
    RECT 27.16 45.48 27.32 46.24 ;
    RECT 27.8 45.48 28.02 46.24 ;
    RECT 28.5 45.48 28.72 46.24 ;
    RECT 29.2 45.48 30.815 46.24 ;
    RECT 31.295 45.48 31.515 46.24 ;
    RECT 31.995 45.48 32.21 46.24 ;
    RECT 32.69 45.48 32.91 46.24 ;
    RECT 33.39 45.48 33.61 46.24 ;
    RECT 34.09 45.48 34.31 46.24 ;
    RECT 34.79 45.48 35.005 46.24 ;
    RECT 35.485 45.48 36.405 46.24 ;
    RECT 36.885 45.48 37.105 46.24 ;
    RECT 37.585 45.48 37.8 46.24 ;
    RECT 38.28 45.48 38.5 46.24 ;
    RECT 38.98 45.48 39.2 46.24 ;
    RECT 39.68 45.48 39.895 46.24 ;
    RECT 40.375 45.48 40.595 46.24 ;
    RECT 41.075 45.48 41.995 46.24 ;
    RECT 42.475 45.48 42.69 46.24 ;
    RECT 43.17 45.48 43.39 46.24 ;
    RECT 43.87 45.48 44.09 46.24 ;
    RECT 44.57 45.48 44.79 46.24 ;
    RECT 45.27 45.48 45.485 46.24 ;
    RECT 45.965 45.48 46.185 46.24 ;
    RECT 46.665 45.48 47.58 46.24 ;
    RECT 48.06 45.48 48.28 46.24 ;
    RECT 48.76 45.48 48.98 46.24 ;
    RECT 49.46 45.48 49.68 46.24 ;
    RECT 50.16 45.48 50.375 46.24 ;
    RECT 50.855 45.48 51.775 46.24 ;
    RECT 52.255 45.48 53.17 46.24 ;
    RECT 53.65 45.48 53.87 46.24 ;
    RECT 54.35 45.48 54.57 46.24 ;
    RECT 55.05 45.48 55.265 46.24 ;
    RECT 55.745 45.48 55.965 46.24 ;
    RECT 56.445 45.48 56.665 46.24 ;
    RECT 57.145 45.48 58.06 46.24 ;
    RECT 58.54 45.48 59.46 46.24 ;
    RECT 59.94 45.48 60.16 46.24 ;
    RECT 60.64 45.48 60.855 46.24 ;
    RECT 61.335 45.48 61.555 46.24 ;
    RECT 62.035 45.48 62.25 46.24 ;
    RECT 62.73 45.48 63.65 46.24 ;
    RECT 64.13 45.48 64.345 46.24 ;
    RECT 64.825 45.48 65.045 46.24 ;
    RECT 65.525 45.48 65.745 46.24 ;
    RECT 66.225 45.48 66.445 46.24 ;
    RECT 66.925 45.48 67.14 46.24 ;
    RECT 67.62 45.48 67.84 46.24 ;
    RECT 68.32 45.48 69.235 46.24 ;
    RECT 69.715 45.48 69.935 46.24 ;
    RECT 70.415 45.48 70.635 46.24 ;
    RECT 71.115 45.48 71.335 46.24 ;
    RECT 71.815 45.48 72.035 46.24 ;
    RECT 72.515 45.48 72.735 46.24 ;
    RECT 73.215 45.48 73.435 46.24 ;
    RECT 73.915 45.48 74.835 46.24 ;
    RECT 75.315 45.48 75.535 46.24 ;
    RECT 76.015 45.48 76.225 46.24 ;
    RECT 76.705 45.48 76.92 46.24 ;
    RECT 77.4 45.48 77.62 46.24 ;
    RECT 78.1 45.48 78.32 46.24 ;
    RECT 78.8 45.48 79.02 46.24 ;
    RECT 79.5 45.48 81.115 46.24 ;
    RECT 81.595 45.48 81.815 46.24 ;
    RECT 82.295 45.48 82.515 46.24 ;
    RECT 82.995 45.48 83.055 46.24 ;
    RECT 83.055 45.39 83.335 46.33 ;
    RECT 83.335 45.48 83.505 46.24 ;
    RECT 26.71 44.72 26.88 45.48 ;
    RECT 26.88 44.63 27.16 45.57 ;
    RECT 27.16 44.72 27.32 45.48 ;
    RECT 27.8 44.72 28.02 45.48 ;
    RECT 28.5 44.72 28.72 45.48 ;
    RECT 29.2 44.72 30.815 45.48 ;
    RECT 31.295 44.72 31.515 45.48 ;
    RECT 31.995 44.72 32.21 45.48 ;
    RECT 32.69 44.72 32.91 45.48 ;
    RECT 33.39 44.72 33.61 45.48 ;
    RECT 34.09 44.72 34.31 45.48 ;
    RECT 34.79 44.72 35.005 45.48 ;
    RECT 35.485 44.72 36.405 45.48 ;
    RECT 36.885 44.72 37.105 45.48 ;
    RECT 37.585 44.72 37.8 45.48 ;
    RECT 38.28 44.72 38.5 45.48 ;
    RECT 38.98 44.72 39.2 45.48 ;
    RECT 39.68 44.72 39.895 45.48 ;
    RECT 40.375 44.72 40.595 45.48 ;
    RECT 41.075 44.72 41.995 45.48 ;
    RECT 42.475 44.72 42.69 45.48 ;
    RECT 43.17 44.72 43.39 45.48 ;
    RECT 43.87 44.72 44.09 45.48 ;
    RECT 44.57 44.72 44.79 45.48 ;
    RECT 45.27 44.72 45.485 45.48 ;
    RECT 45.965 44.72 46.185 45.48 ;
    RECT 46.665 44.72 47.58 45.48 ;
    RECT 48.06 44.72 48.28 45.48 ;
    RECT 48.76 44.72 48.98 45.48 ;
    RECT 49.46 44.72 49.68 45.48 ;
    RECT 50.16 44.72 50.375 45.48 ;
    RECT 50.855 44.72 51.775 45.48 ;
    RECT 52.255 44.72 53.17 45.48 ;
    RECT 53.65 44.72 53.87 45.48 ;
    RECT 54.35 44.72 54.57 45.48 ;
    RECT 55.05 44.72 55.265 45.48 ;
    RECT 55.745 44.72 55.965 45.48 ;
    RECT 56.445 44.72 56.665 45.48 ;
    RECT 57.145 44.72 58.06 45.48 ;
    RECT 58.54 44.72 59.46 45.48 ;
    RECT 59.94 44.72 60.16 45.48 ;
    RECT 60.64 44.72 60.855 45.48 ;
    RECT 61.335 44.72 61.555 45.48 ;
    RECT 62.035 44.72 62.25 45.48 ;
    RECT 62.73 44.72 63.65 45.48 ;
    RECT 64.13 44.72 64.345 45.48 ;
    RECT 64.825 44.72 65.045 45.48 ;
    RECT 65.525 44.72 65.745 45.48 ;
    RECT 66.225 44.72 66.445 45.48 ;
    RECT 66.925 44.72 67.14 45.48 ;
    RECT 67.62 44.72 67.84 45.48 ;
    RECT 68.32 44.72 69.235 45.48 ;
    RECT 69.715 44.72 69.935 45.48 ;
    RECT 70.415 44.72 70.635 45.48 ;
    RECT 71.115 44.72 71.335 45.48 ;
    RECT 71.815 44.72 72.035 45.48 ;
    RECT 72.515 44.72 72.735 45.48 ;
    RECT 73.215 44.72 73.435 45.48 ;
    RECT 73.915 44.72 74.835 45.48 ;
    RECT 75.315 44.72 75.535 45.48 ;
    RECT 76.015 44.72 76.225 45.48 ;
    RECT 76.705 44.72 76.92 45.48 ;
    RECT 77.4 44.72 77.62 45.48 ;
    RECT 78.1 44.72 78.32 45.48 ;
    RECT 78.8 44.72 79.02 45.48 ;
    RECT 79.5 44.72 81.115 45.48 ;
    RECT 81.595 44.72 81.815 45.48 ;
    RECT 82.295 44.72 82.515 45.48 ;
    RECT 82.995 44.72 83.055 45.48 ;
    RECT 83.055 44.63 83.335 45.57 ;
    RECT 83.335 44.72 83.505 45.48 ;
    RECT 26.71 43.96 26.88 44.72 ;
    RECT 26.88 43.87 27.16 44.81 ;
    RECT 27.16 43.96 27.32 44.72 ;
    RECT 27.8 43.96 28.02 44.72 ;
    RECT 28.5 43.96 28.72 44.72 ;
    RECT 29.2 43.96 30.815 44.72 ;
    RECT 31.295 43.96 31.515 44.72 ;
    RECT 31.995 43.96 32.21 44.72 ;
    RECT 32.69 43.96 32.91 44.72 ;
    RECT 33.39 43.96 33.61 44.72 ;
    RECT 34.09 43.96 34.31 44.72 ;
    RECT 34.79 43.96 35.005 44.72 ;
    RECT 35.485 43.96 36.405 44.72 ;
    RECT 36.885 43.96 37.105 44.72 ;
    RECT 37.585 43.96 37.8 44.72 ;
    RECT 38.28 43.96 38.5 44.72 ;
    RECT 38.98 43.96 39.2 44.72 ;
    RECT 39.68 43.96 39.895 44.72 ;
    RECT 40.375 43.96 40.595 44.72 ;
    RECT 41.075 43.96 41.995 44.72 ;
    RECT 42.475 43.96 42.69 44.72 ;
    RECT 43.17 43.96 43.39 44.72 ;
    RECT 43.87 43.96 44.09 44.72 ;
    RECT 44.57 43.96 44.79 44.72 ;
    RECT 45.27 43.96 45.485 44.72 ;
    RECT 45.965 43.96 46.185 44.72 ;
    RECT 46.665 43.96 47.58 44.72 ;
    RECT 48.06 43.96 48.28 44.72 ;
    RECT 48.76 43.96 48.98 44.72 ;
    RECT 49.46 43.96 49.68 44.72 ;
    RECT 50.16 43.96 50.375 44.72 ;
    RECT 50.855 43.96 51.775 44.72 ;
    RECT 52.255 43.96 53.17 44.72 ;
    RECT 53.65 43.96 53.87 44.72 ;
    RECT 54.35 43.96 54.57 44.72 ;
    RECT 55.05 43.96 55.265 44.72 ;
    RECT 55.745 43.96 55.965 44.72 ;
    RECT 56.445 43.96 56.665 44.72 ;
    RECT 57.145 43.96 58.06 44.72 ;
    RECT 58.54 43.96 59.46 44.72 ;
    RECT 59.94 43.96 60.16 44.72 ;
    RECT 60.64 43.96 60.855 44.72 ;
    RECT 61.335 43.96 61.555 44.72 ;
    RECT 62.035 43.96 62.25 44.72 ;
    RECT 62.73 43.96 63.65 44.72 ;
    RECT 64.13 43.96 64.345 44.72 ;
    RECT 64.825 43.96 65.045 44.72 ;
    RECT 65.525 43.96 65.745 44.72 ;
    RECT 66.225 43.96 66.445 44.72 ;
    RECT 66.925 43.96 67.14 44.72 ;
    RECT 67.62 43.96 67.84 44.72 ;
    RECT 68.32 43.96 69.235 44.72 ;
    RECT 69.715 43.96 69.935 44.72 ;
    RECT 70.415 43.96 70.635 44.72 ;
    RECT 71.115 43.96 71.335 44.72 ;
    RECT 71.815 43.96 72.035 44.72 ;
    RECT 72.515 43.96 72.735 44.72 ;
    RECT 73.215 43.96 73.435 44.72 ;
    RECT 73.915 43.96 74.835 44.72 ;
    RECT 75.315 43.96 75.535 44.72 ;
    RECT 76.015 43.96 76.225 44.72 ;
    RECT 76.705 43.96 76.92 44.72 ;
    RECT 77.4 43.96 77.62 44.72 ;
    RECT 78.1 43.96 78.32 44.72 ;
    RECT 78.8 43.96 79.02 44.72 ;
    RECT 79.5 43.96 81.115 44.72 ;
    RECT 81.595 43.96 81.815 44.72 ;
    RECT 82.295 43.96 82.515 44.72 ;
    RECT 82.995 43.96 83.055 44.72 ;
    RECT 83.055 43.87 83.335 44.81 ;
    RECT 83.335 43.96 83.505 44.72 ;
    RECT 26.71 43.2 26.88 43.96 ;
    RECT 26.88 43.11 27.16 44.05 ;
    RECT 27.16 43.2 27.32 43.96 ;
    RECT 27.8 43.2 28.02 43.96 ;
    RECT 28.5 43.2 28.72 43.96 ;
    RECT 29.2 43.2 30.815 43.96 ;
    RECT 31.295 43.2 31.515 43.96 ;
    RECT 31.995 43.2 32.21 43.96 ;
    RECT 32.69 43.2 32.91 43.96 ;
    RECT 33.39 43.2 33.61 43.96 ;
    RECT 34.09 43.2 34.31 43.96 ;
    RECT 34.79 43.2 35.005 43.96 ;
    RECT 35.485 43.2 36.405 43.96 ;
    RECT 36.885 43.2 37.105 43.96 ;
    RECT 37.585 43.2 37.8 43.96 ;
    RECT 38.28 43.2 38.5 43.96 ;
    RECT 38.98 43.2 39.2 43.96 ;
    RECT 39.68 43.2 39.895 43.96 ;
    RECT 40.375 43.2 40.595 43.96 ;
    RECT 41.075 43.2 41.995 43.96 ;
    RECT 42.475 43.2 42.69 43.96 ;
    RECT 43.17 43.2 43.39 43.96 ;
    RECT 43.87 43.2 44.09 43.96 ;
    RECT 44.57 43.2 44.79 43.96 ;
    RECT 45.27 43.2 45.485 43.96 ;
    RECT 45.965 43.2 46.185 43.96 ;
    RECT 46.665 43.2 47.58 43.96 ;
    RECT 48.06 43.2 48.28 43.96 ;
    RECT 48.76 43.2 48.98 43.96 ;
    RECT 49.46 43.2 49.68 43.96 ;
    RECT 50.16 43.2 50.375 43.96 ;
    RECT 50.855 43.2 51.775 43.96 ;
    RECT 52.255 43.2 53.17 43.96 ;
    RECT 53.65 43.2 53.87 43.96 ;
    RECT 54.35 43.2 54.57 43.96 ;
    RECT 55.05 43.2 55.265 43.96 ;
    RECT 55.745 43.2 55.965 43.96 ;
    RECT 56.445 43.2 56.665 43.96 ;
    RECT 57.145 43.2 58.06 43.96 ;
    RECT 58.54 43.2 59.46 43.96 ;
    RECT 59.94 43.2 60.16 43.96 ;
    RECT 60.64 43.2 60.855 43.96 ;
    RECT 61.335 43.2 61.555 43.96 ;
    RECT 62.035 43.2 62.25 43.96 ;
    RECT 62.73 43.2 63.65 43.96 ;
    RECT 64.13 43.2 64.345 43.96 ;
    RECT 64.825 43.2 65.045 43.96 ;
    RECT 65.525 43.2 65.745 43.96 ;
    RECT 66.225 43.2 66.445 43.96 ;
    RECT 66.925 43.2 67.14 43.96 ;
    RECT 67.62 43.2 67.84 43.96 ;
    RECT 68.32 43.2 69.235 43.96 ;
    RECT 69.715 43.2 69.935 43.96 ;
    RECT 70.415 43.2 70.635 43.96 ;
    RECT 71.115 43.2 71.335 43.96 ;
    RECT 71.815 43.2 72.035 43.96 ;
    RECT 72.515 43.2 72.735 43.96 ;
    RECT 73.215 43.2 73.435 43.96 ;
    RECT 73.915 43.2 74.835 43.96 ;
    RECT 75.315 43.2 75.535 43.96 ;
    RECT 76.015 43.2 76.225 43.96 ;
    RECT 76.705 43.2 76.92 43.96 ;
    RECT 77.4 43.2 77.62 43.96 ;
    RECT 78.1 43.2 78.32 43.96 ;
    RECT 78.8 43.2 79.02 43.96 ;
    RECT 79.5 43.2 81.115 43.96 ;
    RECT 81.595 43.2 81.815 43.96 ;
    RECT 82.295 43.2 82.515 43.96 ;
    RECT 82.995 43.2 83.055 43.96 ;
    RECT 83.055 43.11 83.335 44.05 ;
    RECT 83.335 43.2 83.505 43.96 ;
    RECT 26.71 42.44 26.88 43.2 ;
    RECT 26.88 42.35 27.16 43.29 ;
    RECT 27.16 42.44 27.32 43.2 ;
    RECT 27.8 42.44 28.02 43.2 ;
    RECT 28.5 42.44 28.72 43.2 ;
    RECT 29.2 42.44 30.815 43.2 ;
    RECT 31.295 42.44 31.515 43.2 ;
    RECT 31.995 42.44 32.21 43.2 ;
    RECT 32.69 42.44 32.91 43.2 ;
    RECT 33.39 42.44 33.61 43.2 ;
    RECT 34.09 42.44 34.31 43.2 ;
    RECT 34.79 42.44 35.005 43.2 ;
    RECT 35.485 42.44 36.405 43.2 ;
    RECT 36.885 42.44 37.105 43.2 ;
    RECT 37.585 42.44 37.8 43.2 ;
    RECT 38.28 42.44 38.5 43.2 ;
    RECT 38.98 42.44 39.2 43.2 ;
    RECT 39.68 42.44 39.895 43.2 ;
    RECT 40.375 42.44 40.595 43.2 ;
    RECT 41.075 42.44 41.995 43.2 ;
    RECT 42.475 42.44 42.69 43.2 ;
    RECT 43.17 42.44 43.39 43.2 ;
    RECT 43.87 42.44 44.09 43.2 ;
    RECT 44.57 42.44 44.79 43.2 ;
    RECT 45.27 42.44 45.485 43.2 ;
    RECT 45.965 42.44 46.185 43.2 ;
    RECT 46.665 42.44 47.58 43.2 ;
    RECT 48.06 42.44 48.28 43.2 ;
    RECT 48.76 42.44 48.98 43.2 ;
    RECT 49.46 42.44 49.68 43.2 ;
    RECT 50.16 42.44 50.375 43.2 ;
    RECT 50.855 42.44 51.775 43.2 ;
    RECT 52.255 42.44 53.17 43.2 ;
    RECT 53.65 42.44 53.87 43.2 ;
    RECT 54.35 42.44 54.57 43.2 ;
    RECT 55.05 42.44 55.265 43.2 ;
    RECT 55.745 42.44 55.965 43.2 ;
    RECT 56.445 42.44 56.665 43.2 ;
    RECT 57.145 42.44 58.06 43.2 ;
    RECT 58.54 42.44 59.46 43.2 ;
    RECT 59.94 42.44 60.16 43.2 ;
    RECT 60.64 42.44 60.855 43.2 ;
    RECT 61.335 42.44 61.555 43.2 ;
    RECT 62.035 42.44 62.25 43.2 ;
    RECT 62.73 42.44 63.65 43.2 ;
    RECT 64.13 42.44 64.345 43.2 ;
    RECT 64.825 42.44 65.045 43.2 ;
    RECT 65.525 42.44 65.745 43.2 ;
    RECT 66.225 42.44 66.445 43.2 ;
    RECT 66.925 42.44 67.14 43.2 ;
    RECT 67.62 42.44 67.84 43.2 ;
    RECT 68.32 42.44 69.235 43.2 ;
    RECT 69.715 42.44 69.935 43.2 ;
    RECT 70.415 42.44 70.635 43.2 ;
    RECT 71.115 42.44 71.335 43.2 ;
    RECT 71.815 42.44 72.035 43.2 ;
    RECT 72.515 42.44 72.735 43.2 ;
    RECT 73.215 42.44 73.435 43.2 ;
    RECT 73.915 42.44 74.835 43.2 ;
    RECT 75.315 42.44 75.535 43.2 ;
    RECT 76.015 42.44 76.225 43.2 ;
    RECT 76.705 42.44 76.92 43.2 ;
    RECT 77.4 42.44 77.62 43.2 ;
    RECT 78.1 42.44 78.32 43.2 ;
    RECT 78.8 42.44 79.02 43.2 ;
    RECT 79.5 42.44 81.115 43.2 ;
    RECT 81.595 42.44 81.815 43.2 ;
    RECT 82.295 42.44 82.515 43.2 ;
    RECT 82.995 42.44 83.055 43.2 ;
    RECT 83.055 42.35 83.335 43.29 ;
    RECT 83.335 42.44 83.505 43.2 ;
    RECT 26.71 41.68 26.88 42.44 ;
    RECT 26.88 41.59 27.16 42.53 ;
    RECT 27.16 41.68 27.32 42.44 ;
    RECT 27.8 41.68 28.02 42.44 ;
    RECT 28.5 41.68 28.72 42.44 ;
    RECT 29.2 41.68 30.815 42.44 ;
    RECT 31.295 41.68 31.515 42.44 ;
    RECT 31.995 41.68 32.21 42.44 ;
    RECT 32.69 41.68 32.91 42.44 ;
    RECT 33.39 41.68 33.61 42.44 ;
    RECT 34.09 41.68 34.31 42.44 ;
    RECT 34.79 41.68 35.005 42.44 ;
    RECT 35.485 41.68 36.405 42.44 ;
    RECT 36.885 41.68 37.105 42.44 ;
    RECT 37.585 41.68 37.8 42.44 ;
    RECT 38.28 41.68 38.5 42.44 ;
    RECT 38.98 41.68 39.2 42.44 ;
    RECT 39.68 41.68 39.895 42.44 ;
    RECT 40.375 41.68 40.595 42.44 ;
    RECT 41.075 41.68 41.995 42.44 ;
    RECT 42.475 41.68 42.69 42.44 ;
    RECT 43.17 41.68 43.39 42.44 ;
    RECT 43.87 41.68 44.09 42.44 ;
    RECT 44.57 41.68 44.79 42.44 ;
    RECT 45.27 41.68 45.485 42.44 ;
    RECT 45.965 41.68 46.185 42.44 ;
    RECT 46.665 41.68 47.58 42.44 ;
    RECT 48.06 41.68 48.28 42.44 ;
    RECT 48.76 41.68 48.98 42.44 ;
    RECT 49.46 41.68 49.68 42.44 ;
    RECT 50.16 41.68 50.375 42.44 ;
    RECT 50.855 41.68 51.775 42.44 ;
    RECT 52.255 41.68 53.17 42.44 ;
    RECT 53.65 41.68 53.87 42.44 ;
    RECT 54.35 41.68 54.57 42.44 ;
    RECT 55.05 41.68 55.265 42.44 ;
    RECT 55.745 41.68 55.965 42.44 ;
    RECT 56.445 41.68 56.665 42.44 ;
    RECT 57.145 41.68 58.06 42.44 ;
    RECT 58.54 41.68 59.46 42.44 ;
    RECT 59.94 41.68 60.16 42.44 ;
    RECT 60.64 41.68 60.855 42.44 ;
    RECT 61.335 41.68 61.555 42.44 ;
    RECT 62.035 41.68 62.25 42.44 ;
    RECT 62.73 41.68 63.65 42.44 ;
    RECT 64.13 41.68 64.345 42.44 ;
    RECT 64.825 41.68 65.045 42.44 ;
    RECT 65.525 41.68 65.745 42.44 ;
    RECT 66.225 41.68 66.445 42.44 ;
    RECT 66.925 41.68 67.14 42.44 ;
    RECT 67.62 41.68 67.84 42.44 ;
    RECT 68.32 41.68 69.235 42.44 ;
    RECT 69.715 41.68 69.935 42.44 ;
    RECT 70.415 41.68 70.635 42.44 ;
    RECT 71.115 41.68 71.335 42.44 ;
    RECT 71.815 41.68 72.035 42.44 ;
    RECT 72.515 41.68 72.735 42.44 ;
    RECT 73.215 41.68 73.435 42.44 ;
    RECT 73.915 41.68 74.835 42.44 ;
    RECT 75.315 41.68 75.535 42.44 ;
    RECT 76.015 41.68 76.225 42.44 ;
    RECT 76.705 41.68 76.92 42.44 ;
    RECT 77.4 41.68 77.62 42.44 ;
    RECT 78.1 41.68 78.32 42.44 ;
    RECT 78.8 41.68 79.02 42.44 ;
    RECT 79.5 41.68 81.115 42.44 ;
    RECT 81.595 41.68 81.815 42.44 ;
    RECT 82.295 41.68 82.515 42.44 ;
    RECT 82.995 41.68 83.055 42.44 ;
    RECT 83.055 41.59 83.335 42.53 ;
    RECT 83.335 41.68 83.505 42.44 ;
    RECT 26.71 40.92 26.88 41.68 ;
    RECT 26.88 40.83 27.16 41.77 ;
    RECT 27.16 40.92 27.32 41.68 ;
    RECT 27.8 40.92 28.02 41.68 ;
    RECT 28.5 40.92 28.72 41.68 ;
    RECT 29.2 40.92 30.815 41.68 ;
    RECT 31.295 40.92 31.515 41.68 ;
    RECT 31.995 40.92 32.21 41.68 ;
    RECT 32.69 40.92 32.91 41.68 ;
    RECT 33.39 40.92 33.61 41.68 ;
    RECT 34.09 40.92 34.31 41.68 ;
    RECT 34.79 40.92 35.005 41.68 ;
    RECT 35.485 40.92 36.405 41.68 ;
    RECT 36.885 40.92 37.105 41.68 ;
    RECT 37.585 40.92 37.8 41.68 ;
    RECT 38.28 40.92 38.5 41.68 ;
    RECT 38.98 40.92 39.2 41.68 ;
    RECT 39.68 40.92 39.895 41.68 ;
    RECT 40.375 40.92 40.595 41.68 ;
    RECT 41.075 40.92 41.995 41.68 ;
    RECT 42.475 40.92 42.69 41.68 ;
    RECT 43.17 40.92 43.39 41.68 ;
    RECT 43.87 40.92 44.09 41.68 ;
    RECT 44.57 40.92 44.79 41.68 ;
    RECT 45.27 40.92 45.485 41.68 ;
    RECT 45.965 40.92 46.185 41.68 ;
    RECT 46.665 40.92 47.58 41.68 ;
    RECT 48.06 40.92 48.28 41.68 ;
    RECT 48.76 40.92 48.98 41.68 ;
    RECT 49.46 40.92 49.68 41.68 ;
    RECT 50.16 40.92 50.375 41.68 ;
    RECT 50.855 40.92 51.775 41.68 ;
    RECT 52.255 40.92 53.17 41.68 ;
    RECT 53.65 40.92 53.87 41.68 ;
    RECT 54.35 40.92 54.57 41.68 ;
    RECT 55.05 40.92 55.265 41.68 ;
    RECT 55.745 40.92 55.965 41.68 ;
    RECT 56.445 40.92 56.665 41.68 ;
    RECT 57.145 40.92 58.06 41.68 ;
    RECT 58.54 40.92 59.46 41.68 ;
    RECT 59.94 40.92 60.16 41.68 ;
    RECT 60.64 40.92 60.855 41.68 ;
    RECT 61.335 40.92 61.555 41.68 ;
    RECT 62.035 40.92 62.25 41.68 ;
    RECT 62.73 40.92 63.65 41.68 ;
    RECT 64.13 40.92 64.345 41.68 ;
    RECT 64.825 40.92 65.045 41.68 ;
    RECT 65.525 40.92 65.745 41.68 ;
    RECT 66.225 40.92 66.445 41.68 ;
    RECT 66.925 40.92 67.14 41.68 ;
    RECT 67.62 40.92 67.84 41.68 ;
    RECT 68.32 40.92 69.235 41.68 ;
    RECT 69.715 40.92 69.935 41.68 ;
    RECT 70.415 40.92 70.635 41.68 ;
    RECT 71.115 40.92 71.335 41.68 ;
    RECT 71.815 40.92 72.035 41.68 ;
    RECT 72.515 40.92 72.735 41.68 ;
    RECT 73.215 40.92 73.435 41.68 ;
    RECT 73.915 40.92 74.835 41.68 ;
    RECT 75.315 40.92 75.535 41.68 ;
    RECT 76.015 40.92 76.225 41.68 ;
    RECT 76.705 40.92 76.92 41.68 ;
    RECT 77.4 40.92 77.62 41.68 ;
    RECT 78.1 40.92 78.32 41.68 ;
    RECT 78.8 40.92 79.02 41.68 ;
    RECT 79.5 40.92 81.115 41.68 ;
    RECT 81.595 40.92 81.815 41.68 ;
    RECT 82.295 40.92 82.515 41.68 ;
    RECT 82.995 40.92 83.055 41.68 ;
    RECT 83.055 40.83 83.335 41.77 ;
    RECT 83.335 40.92 83.505 41.68 ;
    RECT 26.71 40.16 26.88 40.92 ;
    RECT 26.88 40.07 27.16 41.01 ;
    RECT 27.16 40.16 27.32 40.92 ;
    RECT 27.8 40.16 28.02 40.92 ;
    RECT 28.5 40.16 28.72 40.92 ;
    RECT 29.2 40.16 30.815 40.92 ;
    RECT 31.295 40.16 31.515 40.92 ;
    RECT 31.995 40.16 32.21 40.92 ;
    RECT 32.69 40.16 32.91 40.92 ;
    RECT 33.39 40.16 33.61 40.92 ;
    RECT 34.09 40.16 34.31 40.92 ;
    RECT 34.79 40.16 35.005 40.92 ;
    RECT 35.485 40.16 36.405 40.92 ;
    RECT 36.885 40.16 37.105 40.92 ;
    RECT 37.585 40.16 37.8 40.92 ;
    RECT 38.28 40.16 38.5 40.92 ;
    RECT 38.98 40.16 39.2 40.92 ;
    RECT 39.68 40.16 39.895 40.92 ;
    RECT 40.375 40.16 40.595 40.92 ;
    RECT 41.075 40.16 41.995 40.92 ;
    RECT 42.475 40.16 42.69 40.92 ;
    RECT 43.17 40.16 43.39 40.92 ;
    RECT 43.87 40.16 44.09 40.92 ;
    RECT 44.57 40.16 44.79 40.92 ;
    RECT 45.27 40.16 45.485 40.92 ;
    RECT 45.965 40.16 46.185 40.92 ;
    RECT 46.665 40.16 47.58 40.92 ;
    RECT 48.06 40.16 48.28 40.92 ;
    RECT 48.76 40.16 48.98 40.92 ;
    RECT 49.46 40.16 49.68 40.92 ;
    RECT 50.16 40.16 50.375 40.92 ;
    RECT 50.855 40.16 51.775 40.92 ;
    RECT 52.255 40.16 53.17 40.92 ;
    RECT 53.65 40.16 53.87 40.92 ;
    RECT 54.35 40.16 54.57 40.92 ;
    RECT 55.05 40.16 55.265 40.92 ;
    RECT 55.745 40.16 55.965 40.92 ;
    RECT 56.445 40.16 56.665 40.92 ;
    RECT 57.145 40.16 58.06 40.92 ;
    RECT 58.54 40.16 59.46 40.92 ;
    RECT 59.94 40.16 60.16 40.92 ;
    RECT 60.64 40.16 60.855 40.92 ;
    RECT 61.335 40.16 61.555 40.92 ;
    RECT 62.035 40.16 62.25 40.92 ;
    RECT 62.73 40.16 63.65 40.92 ;
    RECT 64.13 40.16 64.345 40.92 ;
    RECT 64.825 40.16 65.045 40.92 ;
    RECT 65.525 40.16 65.745 40.92 ;
    RECT 66.225 40.16 66.445 40.92 ;
    RECT 66.925 40.16 67.14 40.92 ;
    RECT 67.62 40.16 67.84 40.92 ;
    RECT 68.32 40.16 69.235 40.92 ;
    RECT 69.715 40.16 69.935 40.92 ;
    RECT 70.415 40.16 70.635 40.92 ;
    RECT 71.115 40.16 71.335 40.92 ;
    RECT 71.815 40.16 72.035 40.92 ;
    RECT 72.515 40.16 72.735 40.92 ;
    RECT 73.215 40.16 73.435 40.92 ;
    RECT 73.915 40.16 74.835 40.92 ;
    RECT 75.315 40.16 75.535 40.92 ;
    RECT 76.015 40.16 76.225 40.92 ;
    RECT 76.705 40.16 76.92 40.92 ;
    RECT 77.4 40.16 77.62 40.92 ;
    RECT 78.1 40.16 78.32 40.92 ;
    RECT 78.8 40.16 79.02 40.92 ;
    RECT 79.5 40.16 81.115 40.92 ;
    RECT 81.595 40.16 81.815 40.92 ;
    RECT 82.295 40.16 82.515 40.92 ;
    RECT 82.995 40.16 83.055 40.92 ;
    RECT 83.055 40.07 83.335 41.01 ;
    RECT 83.335 40.16 83.505 40.92 ;
    RECT 26.71 39.4 26.88 40.16 ;
    RECT 26.88 39.31 27.16 40.25 ;
    RECT 27.16 39.4 27.32 40.16 ;
    RECT 27.8 39.4 28.02 40.16 ;
    RECT 28.5 39.4 28.72 40.16 ;
    RECT 29.2 39.4 30.815 40.16 ;
    RECT 31.295 39.4 31.515 40.16 ;
    RECT 31.995 39.4 32.21 40.16 ;
    RECT 32.69 39.4 32.91 40.16 ;
    RECT 33.39 39.4 33.61 40.16 ;
    RECT 34.09 39.4 34.31 40.16 ;
    RECT 34.79 39.4 35.005 40.16 ;
    RECT 35.485 39.4 36.405 40.16 ;
    RECT 36.885 39.4 37.105 40.16 ;
    RECT 37.585 39.4 37.8 40.16 ;
    RECT 38.28 39.4 38.5 40.16 ;
    RECT 38.98 39.4 39.2 40.16 ;
    RECT 39.68 39.4 39.895 40.16 ;
    RECT 40.375 39.4 40.595 40.16 ;
    RECT 41.075 39.4 41.995 40.16 ;
    RECT 42.475 39.4 42.69 40.16 ;
    RECT 43.17 39.4 43.39 40.16 ;
    RECT 43.87 39.4 44.09 40.16 ;
    RECT 44.57 39.4 44.79 40.16 ;
    RECT 45.27 39.4 45.485 40.16 ;
    RECT 45.965 39.4 46.185 40.16 ;
    RECT 46.665 39.4 47.58 40.16 ;
    RECT 48.06 39.4 48.28 40.16 ;
    RECT 48.76 39.4 48.98 40.16 ;
    RECT 49.46 39.4 49.68 40.16 ;
    RECT 50.16 39.4 50.375 40.16 ;
    RECT 50.855 39.4 51.775 40.16 ;
    RECT 52.255 39.4 53.17 40.16 ;
    RECT 53.65 39.4 53.87 40.16 ;
    RECT 54.35 39.4 54.57 40.16 ;
    RECT 55.05 39.4 55.265 40.16 ;
    RECT 55.745 39.4 55.965 40.16 ;
    RECT 56.445 39.4 56.665 40.16 ;
    RECT 57.145 39.4 58.06 40.16 ;
    RECT 58.54 39.4 59.46 40.16 ;
    RECT 59.94 39.4 60.16 40.16 ;
    RECT 60.64 39.4 60.855 40.16 ;
    RECT 61.335 39.4 61.555 40.16 ;
    RECT 62.035 39.4 62.25 40.16 ;
    RECT 62.73 39.4 63.65 40.16 ;
    RECT 64.13 39.4 64.345 40.16 ;
    RECT 64.825 39.4 65.045 40.16 ;
    RECT 65.525 39.4 65.745 40.16 ;
    RECT 66.225 39.4 66.445 40.16 ;
    RECT 66.925 39.4 67.14 40.16 ;
    RECT 67.62 39.4 67.84 40.16 ;
    RECT 68.32 39.4 69.235 40.16 ;
    RECT 69.715 39.4 69.935 40.16 ;
    RECT 70.415 39.4 70.635 40.16 ;
    RECT 71.115 39.4 71.335 40.16 ;
    RECT 71.815 39.4 72.035 40.16 ;
    RECT 72.515 39.4 72.735 40.16 ;
    RECT 73.215 39.4 73.435 40.16 ;
    RECT 73.915 39.4 74.835 40.16 ;
    RECT 75.315 39.4 75.535 40.16 ;
    RECT 76.015 39.4 76.225 40.16 ;
    RECT 76.705 39.4 76.92 40.16 ;
    RECT 77.4 39.4 77.62 40.16 ;
    RECT 78.1 39.4 78.32 40.16 ;
    RECT 78.8 39.4 79.02 40.16 ;
    RECT 79.5 39.4 81.115 40.16 ;
    RECT 81.595 39.4 81.815 40.16 ;
    RECT 82.295 39.4 82.515 40.16 ;
    RECT 82.995 39.4 83.055 40.16 ;
    RECT 83.055 39.31 83.335 40.25 ;
    RECT 83.335 39.4 83.505 40.16 ;
    RECT 26.71 38.64 26.88 39.4 ;
    RECT 26.88 38.55 27.16 39.49 ;
    RECT 27.16 38.64 27.32 39.4 ;
    RECT 27.8 38.64 28.02 39.4 ;
    RECT 28.5 38.64 28.72 39.4 ;
    RECT 29.2 38.64 30.815 39.4 ;
    RECT 31.295 38.64 31.515 39.4 ;
    RECT 31.995 38.64 32.21 39.4 ;
    RECT 32.69 38.64 32.91 39.4 ;
    RECT 33.39 38.64 33.61 39.4 ;
    RECT 34.09 38.64 34.31 39.4 ;
    RECT 34.79 38.64 35.005 39.4 ;
    RECT 35.485 38.64 36.405 39.4 ;
    RECT 36.885 38.64 37.105 39.4 ;
    RECT 37.585 38.64 37.8 39.4 ;
    RECT 38.28 38.64 38.5 39.4 ;
    RECT 38.98 38.64 39.2 39.4 ;
    RECT 39.68 38.64 39.895 39.4 ;
    RECT 40.375 38.64 40.595 39.4 ;
    RECT 41.075 38.64 41.995 39.4 ;
    RECT 42.475 38.64 42.69 39.4 ;
    RECT 43.17 38.64 43.39 39.4 ;
    RECT 43.87 38.64 44.09 39.4 ;
    RECT 44.57 38.64 44.79 39.4 ;
    RECT 45.27 38.64 45.485 39.4 ;
    RECT 45.965 38.64 46.185 39.4 ;
    RECT 46.665 38.64 47.58 39.4 ;
    RECT 48.06 38.64 48.28 39.4 ;
    RECT 48.76 38.64 48.98 39.4 ;
    RECT 49.46 38.64 49.68 39.4 ;
    RECT 50.16 38.64 50.375 39.4 ;
    RECT 50.855 38.64 51.775 39.4 ;
    RECT 52.255 38.64 53.17 39.4 ;
    RECT 53.65 38.64 53.87 39.4 ;
    RECT 54.35 38.64 54.57 39.4 ;
    RECT 55.05 38.64 55.265 39.4 ;
    RECT 55.745 38.64 55.965 39.4 ;
    RECT 56.445 38.64 56.665 39.4 ;
    RECT 57.145 38.64 58.06 39.4 ;
    RECT 58.54 38.64 59.46 39.4 ;
    RECT 59.94 38.64 60.16 39.4 ;
    RECT 60.64 38.64 60.855 39.4 ;
    RECT 61.335 38.64 61.555 39.4 ;
    RECT 62.035 38.64 62.25 39.4 ;
    RECT 62.73 38.64 63.65 39.4 ;
    RECT 64.13 38.64 64.345 39.4 ;
    RECT 64.825 38.64 65.045 39.4 ;
    RECT 65.525 38.64 65.745 39.4 ;
    RECT 66.225 38.64 66.445 39.4 ;
    RECT 66.925 38.64 67.14 39.4 ;
    RECT 67.62 38.64 67.84 39.4 ;
    RECT 68.32 38.64 69.235 39.4 ;
    RECT 69.715 38.64 69.935 39.4 ;
    RECT 70.415 38.64 70.635 39.4 ;
    RECT 71.115 38.64 71.335 39.4 ;
    RECT 71.815 38.64 72.035 39.4 ;
    RECT 72.515 38.64 72.735 39.4 ;
    RECT 73.215 38.64 73.435 39.4 ;
    RECT 73.915 38.64 74.835 39.4 ;
    RECT 75.315 38.64 75.535 39.4 ;
    RECT 76.015 38.64 76.225 39.4 ;
    RECT 76.705 38.64 76.92 39.4 ;
    RECT 77.4 38.64 77.62 39.4 ;
    RECT 78.1 38.64 78.32 39.4 ;
    RECT 78.8 38.64 79.02 39.4 ;
    RECT 79.5 38.64 81.115 39.4 ;
    RECT 81.595 38.64 81.815 39.4 ;
    RECT 82.295 38.64 82.515 39.4 ;
    RECT 82.995 38.64 83.055 39.4 ;
    RECT 83.055 38.55 83.335 39.49 ;
    RECT 83.335 38.64 83.505 39.4 ;
    RECT 26.71 37.88 26.88 38.64 ;
    RECT 26.88 37.79 27.16 38.73 ;
    RECT 27.16 37.88 27.32 38.64 ;
    RECT 27.8 37.88 28.02 38.64 ;
    RECT 28.5 37.88 28.72 38.64 ;
    RECT 29.2 37.88 30.815 38.64 ;
    RECT 31.295 37.88 31.515 38.64 ;
    RECT 31.995 37.88 32.21 38.64 ;
    RECT 32.69 37.88 32.91 38.64 ;
    RECT 33.39 37.88 33.61 38.64 ;
    RECT 34.09 37.88 34.31 38.64 ;
    RECT 34.79 37.88 35.005 38.64 ;
    RECT 35.485 37.88 36.405 38.64 ;
    RECT 36.885 37.88 37.105 38.64 ;
    RECT 37.585 37.88 37.8 38.64 ;
    RECT 38.28 37.88 38.5 38.64 ;
    RECT 38.98 37.88 39.2 38.64 ;
    RECT 39.68 37.88 39.895 38.64 ;
    RECT 40.375 37.88 40.595 38.64 ;
    RECT 41.075 37.88 41.995 38.64 ;
    RECT 42.475 37.88 42.69 38.64 ;
    RECT 43.17 37.88 43.39 38.64 ;
    RECT 43.87 37.88 44.09 38.64 ;
    RECT 44.57 37.88 44.79 38.64 ;
    RECT 45.27 37.88 45.485 38.64 ;
    RECT 45.965 37.88 46.185 38.64 ;
    RECT 46.665 37.88 47.58 38.64 ;
    RECT 48.06 37.88 48.28 38.64 ;
    RECT 48.76 37.88 48.98 38.64 ;
    RECT 49.46 37.88 49.68 38.64 ;
    RECT 50.16 37.88 50.375 38.64 ;
    RECT 50.855 37.88 51.775 38.64 ;
    RECT 52.255 37.88 53.17 38.64 ;
    RECT 53.65 37.88 53.87 38.64 ;
    RECT 54.35 37.88 54.57 38.64 ;
    RECT 55.05 37.88 55.265 38.64 ;
    RECT 55.745 37.88 55.965 38.64 ;
    RECT 56.445 37.88 56.665 38.64 ;
    RECT 57.145 37.88 58.06 38.64 ;
    RECT 58.54 37.88 59.46 38.64 ;
    RECT 59.94 37.88 60.16 38.64 ;
    RECT 60.64 37.88 60.855 38.64 ;
    RECT 61.335 37.88 61.555 38.64 ;
    RECT 62.035 37.88 62.25 38.64 ;
    RECT 62.73 37.88 63.65 38.64 ;
    RECT 64.13 37.88 64.345 38.64 ;
    RECT 64.825 37.88 65.045 38.64 ;
    RECT 65.525 37.88 65.745 38.64 ;
    RECT 66.225 37.88 66.445 38.64 ;
    RECT 66.925 37.88 67.14 38.64 ;
    RECT 67.62 37.88 67.84 38.64 ;
    RECT 68.32 37.88 69.235 38.64 ;
    RECT 69.715 37.88 69.935 38.64 ;
    RECT 70.415 37.88 70.635 38.64 ;
    RECT 71.115 37.88 71.335 38.64 ;
    RECT 71.815 37.88 72.035 38.64 ;
    RECT 72.515 37.88 72.735 38.64 ;
    RECT 73.215 37.88 73.435 38.64 ;
    RECT 73.915 37.88 74.835 38.64 ;
    RECT 75.315 37.88 75.535 38.64 ;
    RECT 76.015 37.88 76.225 38.64 ;
    RECT 76.705 37.88 76.92 38.64 ;
    RECT 77.4 37.88 77.62 38.64 ;
    RECT 78.1 37.88 78.32 38.64 ;
    RECT 78.8 37.88 79.02 38.64 ;
    RECT 79.5 37.88 81.115 38.64 ;
    RECT 81.595 37.88 81.815 38.64 ;
    RECT 82.295 37.88 82.515 38.64 ;
    RECT 82.995 37.88 83.055 38.64 ;
    RECT 83.055 37.79 83.335 38.73 ;
    RECT 83.335 37.88 83.505 38.64 ;
    RECT 26.71 37.12 26.88 37.88 ;
    RECT 26.88 37.03 27.16 37.97 ;
    RECT 27.16 37.12 27.32 37.88 ;
    RECT 27.8 37.12 28.02 37.88 ;
    RECT 28.5 37.12 28.72 37.88 ;
    RECT 29.2 37.12 30.815 37.88 ;
    RECT 31.295 37.12 31.515 37.88 ;
    RECT 31.995 37.12 32.21 37.88 ;
    RECT 32.69 37.12 32.91 37.88 ;
    RECT 33.39 37.12 33.61 37.88 ;
    RECT 34.09 37.12 34.31 37.88 ;
    RECT 34.79 37.12 35.005 37.88 ;
    RECT 35.485 37.12 36.405 37.88 ;
    RECT 36.885 37.12 37.105 37.88 ;
    RECT 37.585 37.12 37.8 37.88 ;
    RECT 38.28 37.12 38.5 37.88 ;
    RECT 38.98 37.12 39.2 37.88 ;
    RECT 39.68 37.12 39.895 37.88 ;
    RECT 40.375 37.12 40.595 37.88 ;
    RECT 41.075 37.12 41.995 37.88 ;
    RECT 42.475 37.12 42.69 37.88 ;
    RECT 43.17 37.12 43.39 37.88 ;
    RECT 43.87 37.12 44.09 37.88 ;
    RECT 44.57 37.12 44.79 37.88 ;
    RECT 45.27 37.12 45.485 37.88 ;
    RECT 45.965 37.12 46.185 37.88 ;
    RECT 46.665 37.12 47.58 37.88 ;
    RECT 48.06 37.12 48.28 37.88 ;
    RECT 48.76 37.12 48.98 37.88 ;
    RECT 49.46 37.12 49.68 37.88 ;
    RECT 50.16 37.12 50.375 37.88 ;
    RECT 50.855 37.12 51.775 37.88 ;
    RECT 52.255 37.12 53.17 37.88 ;
    RECT 53.65 37.12 53.87 37.88 ;
    RECT 54.35 37.12 54.57 37.88 ;
    RECT 55.05 37.12 55.265 37.88 ;
    RECT 55.745 37.12 55.965 37.88 ;
    RECT 56.445 37.12 56.665 37.88 ;
    RECT 57.145 37.12 58.06 37.88 ;
    RECT 58.54 37.12 59.46 37.88 ;
    RECT 59.94 37.12 60.16 37.88 ;
    RECT 60.64 37.12 60.855 37.88 ;
    RECT 61.335 37.12 61.555 37.88 ;
    RECT 62.035 37.12 62.25 37.88 ;
    RECT 62.73 37.12 63.65 37.88 ;
    RECT 64.13 37.12 64.345 37.88 ;
    RECT 64.825 37.12 65.045 37.88 ;
    RECT 65.525 37.12 65.745 37.88 ;
    RECT 66.225 37.12 66.445 37.88 ;
    RECT 66.925 37.12 67.14 37.88 ;
    RECT 67.62 37.12 67.84 37.88 ;
    RECT 68.32 37.12 69.235 37.88 ;
    RECT 69.715 37.12 69.935 37.88 ;
    RECT 70.415 37.12 70.635 37.88 ;
    RECT 71.115 37.12 71.335 37.88 ;
    RECT 71.815 37.12 72.035 37.88 ;
    RECT 72.515 37.12 72.735 37.88 ;
    RECT 73.215 37.12 73.435 37.88 ;
    RECT 73.915 37.12 74.835 37.88 ;
    RECT 75.315 37.12 75.535 37.88 ;
    RECT 76.015 37.12 76.225 37.88 ;
    RECT 76.705 37.12 76.92 37.88 ;
    RECT 77.4 37.12 77.62 37.88 ;
    RECT 78.1 37.12 78.32 37.88 ;
    RECT 78.8 37.12 79.02 37.88 ;
    RECT 79.5 37.12 81.115 37.88 ;
    RECT 81.595 37.12 81.815 37.88 ;
    RECT 82.295 37.12 82.515 37.88 ;
    RECT 82.995 37.12 83.055 37.88 ;
    RECT 83.055 37.03 83.335 37.97 ;
    RECT 83.335 37.12 83.505 37.88 ;
    RECT 26.71 36.36 26.88 37.12 ;
    RECT 26.88 36.27 27.16 37.21 ;
    RECT 27.16 36.36 27.32 37.12 ;
    RECT 27.8 36.36 28.02 37.12 ;
    RECT 28.5 36.36 28.72 37.12 ;
    RECT 29.2 36.36 30.815 37.12 ;
    RECT 31.295 36.36 31.515 37.12 ;
    RECT 31.995 36.36 32.21 37.12 ;
    RECT 32.69 36.36 32.91 37.12 ;
    RECT 33.39 36.36 33.61 37.12 ;
    RECT 34.09 36.36 34.31 37.12 ;
    RECT 34.79 36.36 35.005 37.12 ;
    RECT 35.485 36.36 36.405 37.12 ;
    RECT 36.885 36.36 37.105 37.12 ;
    RECT 37.585 36.36 37.8 37.12 ;
    RECT 38.28 36.36 38.5 37.12 ;
    RECT 38.98 36.36 39.2 37.12 ;
    RECT 39.68 36.36 39.895 37.12 ;
    RECT 40.375 36.36 40.595 37.12 ;
    RECT 41.075 36.36 41.995 37.12 ;
    RECT 42.475 36.36 42.69 37.12 ;
    RECT 43.17 36.36 43.39 37.12 ;
    RECT 43.87 36.36 44.09 37.12 ;
    RECT 44.57 36.36 44.79 37.12 ;
    RECT 45.27 36.36 45.485 37.12 ;
    RECT 45.965 36.36 46.185 37.12 ;
    RECT 46.665 36.36 47.58 37.12 ;
    RECT 48.06 36.36 48.28 37.12 ;
    RECT 48.76 36.36 48.98 37.12 ;
    RECT 49.46 36.36 49.68 37.12 ;
    RECT 50.16 36.36 50.375 37.12 ;
    RECT 50.855 36.36 51.775 37.12 ;
    RECT 52.255 36.36 53.17 37.12 ;
    RECT 53.65 36.36 53.87 37.12 ;
    RECT 54.35 36.36 54.57 37.12 ;
    RECT 55.05 36.36 55.265 37.12 ;
    RECT 55.745 36.36 55.965 37.12 ;
    RECT 56.445 36.36 56.665 37.12 ;
    RECT 57.145 36.36 58.06 37.12 ;
    RECT 58.54 36.36 59.46 37.12 ;
    RECT 59.94 36.36 60.16 37.12 ;
    RECT 60.64 36.36 60.855 37.12 ;
    RECT 61.335 36.36 61.555 37.12 ;
    RECT 62.035 36.36 62.25 37.12 ;
    RECT 62.73 36.36 63.65 37.12 ;
    RECT 64.13 36.36 64.345 37.12 ;
    RECT 64.825 36.36 65.045 37.12 ;
    RECT 65.525 36.36 65.745 37.12 ;
    RECT 66.225 36.36 66.445 37.12 ;
    RECT 66.925 36.36 67.14 37.12 ;
    RECT 67.62 36.36 67.84 37.12 ;
    RECT 68.32 36.36 69.235 37.12 ;
    RECT 69.715 36.36 69.935 37.12 ;
    RECT 70.415 36.36 70.635 37.12 ;
    RECT 71.115 36.36 71.335 37.12 ;
    RECT 71.815 36.36 72.035 37.12 ;
    RECT 72.515 36.36 72.735 37.12 ;
    RECT 73.215 36.36 73.435 37.12 ;
    RECT 73.915 36.36 74.835 37.12 ;
    RECT 75.315 36.36 75.535 37.12 ;
    RECT 76.015 36.36 76.225 37.12 ;
    RECT 76.705 36.36 76.92 37.12 ;
    RECT 77.4 36.36 77.62 37.12 ;
    RECT 78.1 36.36 78.32 37.12 ;
    RECT 78.8 36.36 79.02 37.12 ;
    RECT 79.5 36.36 81.115 37.12 ;
    RECT 81.595 36.36 81.815 37.12 ;
    RECT 82.295 36.36 82.515 37.12 ;
    RECT 82.995 36.36 83.055 37.12 ;
    RECT 83.055 36.27 83.335 37.21 ;
    RECT 83.335 36.36 83.505 37.12 ;
    RECT 26.71 35.6 26.88 36.36 ;
    RECT 26.88 35.51 27.16 36.45 ;
    RECT 27.16 35.6 27.32 36.36 ;
    RECT 27.8 35.6 28.02 36.36 ;
    RECT 28.5 35.6 28.72 36.36 ;
    RECT 29.2 35.6 30.815 36.36 ;
    RECT 31.295 35.6 31.515 36.36 ;
    RECT 31.995 35.6 32.21 36.36 ;
    RECT 32.69 35.6 32.91 36.36 ;
    RECT 33.39 35.6 33.61 36.36 ;
    RECT 34.09 35.6 34.31 36.36 ;
    RECT 34.79 35.6 35.005 36.36 ;
    RECT 35.485 35.6 36.405 36.36 ;
    RECT 36.885 35.6 37.105 36.36 ;
    RECT 37.585 35.6 37.8 36.36 ;
    RECT 38.28 35.6 38.5 36.36 ;
    RECT 38.98 35.6 39.2 36.36 ;
    RECT 39.68 35.6 39.895 36.36 ;
    RECT 40.375 35.6 40.595 36.36 ;
    RECT 41.075 35.6 41.995 36.36 ;
    RECT 42.475 35.6 42.69 36.36 ;
    RECT 43.17 35.6 43.39 36.36 ;
    RECT 43.87 35.6 44.09 36.36 ;
    RECT 44.57 35.6 44.79 36.36 ;
    RECT 45.27 35.6 45.485 36.36 ;
    RECT 45.965 35.6 46.185 36.36 ;
    RECT 46.665 35.6 47.58 36.36 ;
    RECT 48.06 35.6 48.28 36.36 ;
    RECT 48.76 35.6 48.98 36.36 ;
    RECT 49.46 35.6 49.68 36.36 ;
    RECT 50.16 35.6 50.375 36.36 ;
    RECT 50.855 35.6 51.775 36.36 ;
    RECT 52.255 35.6 53.17 36.36 ;
    RECT 53.65 35.6 53.87 36.36 ;
    RECT 54.35 35.6 54.57 36.36 ;
    RECT 55.05 35.6 55.265 36.36 ;
    RECT 55.745 35.6 55.965 36.36 ;
    RECT 56.445 35.6 56.665 36.36 ;
    RECT 57.145 35.6 58.06 36.36 ;
    RECT 58.54 35.6 59.46 36.36 ;
    RECT 59.94 35.6 60.16 36.36 ;
    RECT 60.64 35.6 60.855 36.36 ;
    RECT 61.335 35.6 61.555 36.36 ;
    RECT 62.035 35.6 62.25 36.36 ;
    RECT 62.73 35.6 63.65 36.36 ;
    RECT 64.13 35.6 64.345 36.36 ;
    RECT 64.825 35.6 65.045 36.36 ;
    RECT 65.525 35.6 65.745 36.36 ;
    RECT 66.225 35.6 66.445 36.36 ;
    RECT 66.925 35.6 67.14 36.36 ;
    RECT 67.62 35.6 67.84 36.36 ;
    RECT 68.32 35.6 69.235 36.36 ;
    RECT 69.715 35.6 69.935 36.36 ;
    RECT 70.415 35.6 70.635 36.36 ;
    RECT 71.115 35.6 71.335 36.36 ;
    RECT 71.815 35.6 72.035 36.36 ;
    RECT 72.515 35.6 72.735 36.36 ;
    RECT 73.215 35.6 73.435 36.36 ;
    RECT 73.915 35.6 74.835 36.36 ;
    RECT 75.315 35.6 75.535 36.36 ;
    RECT 76.015 35.6 76.225 36.36 ;
    RECT 76.705 35.6 76.92 36.36 ;
    RECT 77.4 35.6 77.62 36.36 ;
    RECT 78.1 35.6 78.32 36.36 ;
    RECT 78.8 35.6 79.02 36.36 ;
    RECT 79.5 35.6 81.115 36.36 ;
    RECT 81.595 35.6 81.815 36.36 ;
    RECT 82.295 35.6 82.515 36.36 ;
    RECT 82.995 35.6 83.055 36.36 ;
    RECT 83.055 35.51 83.335 36.45 ;
    RECT 83.335 35.6 83.505 36.36 ;
    RECT 26.71 34.84 26.88 35.6 ;
    RECT 26.88 34.75 27.16 35.69 ;
    RECT 27.16 34.84 27.32 35.6 ;
    RECT 27.8 34.84 28.02 35.6 ;
    RECT 28.5 34.84 28.72 35.6 ;
    RECT 29.2 34.84 30.815 35.6 ;
    RECT 31.295 34.84 31.515 35.6 ;
    RECT 31.995 34.84 32.21 35.6 ;
    RECT 32.69 34.84 32.91 35.6 ;
    RECT 33.39 34.84 33.61 35.6 ;
    RECT 34.09 34.84 34.31 35.6 ;
    RECT 34.79 34.84 35.005 35.6 ;
    RECT 35.485 34.84 36.405 35.6 ;
    RECT 36.885 34.84 37.105 35.6 ;
    RECT 37.585 34.84 37.8 35.6 ;
    RECT 38.28 34.84 38.5 35.6 ;
    RECT 38.98 34.84 39.2 35.6 ;
    RECT 39.68 34.84 39.895 35.6 ;
    RECT 40.375 34.84 40.595 35.6 ;
    RECT 41.075 34.84 41.995 35.6 ;
    RECT 42.475 34.84 42.69 35.6 ;
    RECT 43.17 34.84 43.39 35.6 ;
    RECT 43.87 34.84 44.09 35.6 ;
    RECT 44.57 34.84 44.79 35.6 ;
    RECT 45.27 34.84 45.485 35.6 ;
    RECT 45.965 34.84 46.185 35.6 ;
    RECT 46.665 34.84 47.58 35.6 ;
    RECT 48.06 34.84 48.28 35.6 ;
    RECT 48.76 34.84 48.98 35.6 ;
    RECT 49.46 34.84 49.68 35.6 ;
    RECT 50.16 34.84 50.375 35.6 ;
    RECT 50.855 34.84 51.775 35.6 ;
    RECT 52.255 34.84 53.17 35.6 ;
    RECT 53.65 34.84 53.87 35.6 ;
    RECT 54.35 34.84 54.57 35.6 ;
    RECT 55.05 34.84 55.265 35.6 ;
    RECT 55.745 34.84 55.965 35.6 ;
    RECT 56.445 34.84 56.665 35.6 ;
    RECT 57.145 34.84 58.06 35.6 ;
    RECT 58.54 34.84 59.46 35.6 ;
    RECT 59.94 34.84 60.16 35.6 ;
    RECT 60.64 34.84 60.855 35.6 ;
    RECT 61.335 34.84 61.555 35.6 ;
    RECT 62.035 34.84 62.25 35.6 ;
    RECT 62.73 34.84 63.65 35.6 ;
    RECT 64.13 34.84 64.345 35.6 ;
    RECT 64.825 34.84 65.045 35.6 ;
    RECT 65.525 34.84 65.745 35.6 ;
    RECT 66.225 34.84 66.445 35.6 ;
    RECT 66.925 34.84 67.14 35.6 ;
    RECT 67.62 34.84 67.84 35.6 ;
    RECT 68.32 34.84 69.235 35.6 ;
    RECT 69.715 34.84 69.935 35.6 ;
    RECT 70.415 34.84 70.635 35.6 ;
    RECT 71.115 34.84 71.335 35.6 ;
    RECT 71.815 34.84 72.035 35.6 ;
    RECT 72.515 34.84 72.735 35.6 ;
    RECT 73.215 34.84 73.435 35.6 ;
    RECT 73.915 34.84 74.835 35.6 ;
    RECT 75.315 34.84 75.535 35.6 ;
    RECT 76.015 34.84 76.225 35.6 ;
    RECT 76.705 34.84 76.92 35.6 ;
    RECT 77.4 34.84 77.62 35.6 ;
    RECT 78.1 34.84 78.32 35.6 ;
    RECT 78.8 34.84 79.02 35.6 ;
    RECT 79.5 34.84 81.115 35.6 ;
    RECT 81.595 34.84 81.815 35.6 ;
    RECT 82.295 34.84 82.515 35.6 ;
    RECT 82.995 34.84 83.055 35.6 ;
    RECT 83.055 34.75 83.335 35.69 ;
    RECT 83.335 34.84 83.505 35.6 ;
    RECT 26.71 34.08 26.88 34.84 ;
    RECT 26.88 33.99 27.16 34.93 ;
    RECT 27.16 34.08 27.32 34.84 ;
    RECT 27.8 34.08 28.02 34.84 ;
    RECT 28.5 34.08 28.72 34.84 ;
    RECT 29.2 34.08 30.815 34.84 ;
    RECT 31.295 34.08 31.515 34.84 ;
    RECT 31.995 34.08 32.21 34.84 ;
    RECT 32.69 34.08 32.91 34.84 ;
    RECT 33.39 34.08 33.61 34.84 ;
    RECT 34.09 34.08 34.31 34.84 ;
    RECT 34.79 34.08 35.005 34.84 ;
    RECT 35.485 34.08 36.405 34.84 ;
    RECT 36.885 34.08 37.105 34.84 ;
    RECT 37.585 34.08 37.8 34.84 ;
    RECT 38.28 34.08 38.5 34.84 ;
    RECT 38.98 34.08 39.2 34.84 ;
    RECT 39.68 34.08 39.895 34.84 ;
    RECT 40.375 34.08 40.595 34.84 ;
    RECT 41.075 34.08 41.995 34.84 ;
    RECT 42.475 34.08 42.69 34.84 ;
    RECT 43.17 34.08 43.39 34.84 ;
    RECT 43.87 34.08 44.09 34.84 ;
    RECT 44.57 34.08 44.79 34.84 ;
    RECT 45.27 34.08 45.485 34.84 ;
    RECT 45.965 34.08 46.185 34.84 ;
    RECT 46.665 34.08 47.58 34.84 ;
    RECT 48.06 34.08 48.28 34.84 ;
    RECT 48.76 34.08 48.98 34.84 ;
    RECT 49.46 34.08 49.68 34.84 ;
    RECT 50.16 34.08 50.375 34.84 ;
    RECT 50.855 34.08 51.775 34.84 ;
    RECT 52.255 34.08 53.17 34.84 ;
    RECT 53.65 34.08 53.87 34.84 ;
    RECT 54.35 34.08 54.57 34.84 ;
    RECT 55.05 34.08 55.265 34.84 ;
    RECT 55.745 34.08 55.965 34.84 ;
    RECT 56.445 34.08 56.665 34.84 ;
    RECT 57.145 34.08 58.06 34.84 ;
    RECT 58.54 34.08 59.46 34.84 ;
    RECT 59.94 34.08 60.16 34.84 ;
    RECT 60.64 34.08 60.855 34.84 ;
    RECT 61.335 34.08 61.555 34.84 ;
    RECT 62.035 34.08 62.25 34.84 ;
    RECT 62.73 34.08 63.65 34.84 ;
    RECT 64.13 34.08 64.345 34.84 ;
    RECT 64.825 34.08 65.045 34.84 ;
    RECT 65.525 34.08 65.745 34.84 ;
    RECT 66.225 34.08 66.445 34.84 ;
    RECT 66.925 34.08 67.14 34.84 ;
    RECT 67.62 34.08 67.84 34.84 ;
    RECT 68.32 34.08 69.235 34.84 ;
    RECT 69.715 34.08 69.935 34.84 ;
    RECT 70.415 34.08 70.635 34.84 ;
    RECT 71.115 34.08 71.335 34.84 ;
    RECT 71.815 34.08 72.035 34.84 ;
    RECT 72.515 34.08 72.735 34.84 ;
    RECT 73.215 34.08 73.435 34.84 ;
    RECT 73.915 34.08 74.835 34.84 ;
    RECT 75.315 34.08 75.535 34.84 ;
    RECT 76.015 34.08 76.225 34.84 ;
    RECT 76.705 34.08 76.92 34.84 ;
    RECT 77.4 34.08 77.62 34.84 ;
    RECT 78.1 34.08 78.32 34.84 ;
    RECT 78.8 34.08 79.02 34.84 ;
    RECT 79.5 34.08 81.115 34.84 ;
    RECT 81.595 34.08 81.815 34.84 ;
    RECT 82.295 34.08 82.515 34.84 ;
    RECT 82.995 34.08 83.055 34.84 ;
    RECT 83.055 33.99 83.335 34.93 ;
    RECT 83.335 34.08 83.505 34.84 ;
    RECT 26.71 33.32 26.88 34.08 ;
    RECT 26.88 33.23 27.16 34.17 ;
    RECT 27.16 33.32 27.32 34.08 ;
    RECT 27.8 33.32 28.02 34.08 ;
    RECT 28.5 33.32 28.72 34.08 ;
    RECT 29.2 33.32 30.815 34.08 ;
    RECT 31.295 33.32 31.515 34.08 ;
    RECT 31.995 33.32 32.21 34.08 ;
    RECT 32.69 33.32 32.91 34.08 ;
    RECT 33.39 33.32 33.61 34.08 ;
    RECT 34.09 33.32 34.31 34.08 ;
    RECT 34.79 33.32 35.005 34.08 ;
    RECT 35.485 33.32 36.405 34.08 ;
    RECT 36.885 33.32 37.105 34.08 ;
    RECT 37.585 33.32 37.8 34.08 ;
    RECT 38.28 33.32 38.5 34.08 ;
    RECT 38.98 33.32 39.2 34.08 ;
    RECT 39.68 33.32 39.895 34.08 ;
    RECT 40.375 33.32 40.595 34.08 ;
    RECT 41.075 33.32 41.995 34.08 ;
    RECT 42.475 33.32 42.69 34.08 ;
    RECT 43.17 33.32 43.39 34.08 ;
    RECT 43.87 33.32 44.09 34.08 ;
    RECT 44.57 33.32 44.79 34.08 ;
    RECT 45.27 33.32 45.485 34.08 ;
    RECT 45.965 33.32 46.185 34.08 ;
    RECT 46.665 33.32 47.58 34.08 ;
    RECT 48.06 33.32 48.28 34.08 ;
    RECT 48.76 33.32 48.98 34.08 ;
    RECT 49.46 33.32 49.68 34.08 ;
    RECT 50.16 33.32 50.375 34.08 ;
    RECT 50.855 33.32 51.775 34.08 ;
    RECT 52.255 33.32 53.17 34.08 ;
    RECT 53.65 33.32 53.87 34.08 ;
    RECT 54.35 33.32 54.57 34.08 ;
    RECT 55.05 33.32 55.265 34.08 ;
    RECT 55.745 33.32 55.965 34.08 ;
    RECT 56.445 33.32 56.665 34.08 ;
    RECT 57.145 33.32 58.06 34.08 ;
    RECT 58.54 33.32 59.46 34.08 ;
    RECT 59.94 33.32 60.16 34.08 ;
    RECT 60.64 33.32 60.855 34.08 ;
    RECT 61.335 33.32 61.555 34.08 ;
    RECT 62.035 33.32 62.25 34.08 ;
    RECT 62.73 33.32 63.65 34.08 ;
    RECT 64.13 33.32 64.345 34.08 ;
    RECT 64.825 33.32 65.045 34.08 ;
    RECT 65.525 33.32 65.745 34.08 ;
    RECT 66.225 33.32 66.445 34.08 ;
    RECT 66.925 33.32 67.14 34.08 ;
    RECT 67.62 33.32 67.84 34.08 ;
    RECT 68.32 33.32 69.235 34.08 ;
    RECT 69.715 33.32 69.935 34.08 ;
    RECT 70.415 33.32 70.635 34.08 ;
    RECT 71.115 33.32 71.335 34.08 ;
    RECT 71.815 33.32 72.035 34.08 ;
    RECT 72.515 33.32 72.735 34.08 ;
    RECT 73.215 33.32 73.435 34.08 ;
    RECT 73.915 33.32 74.835 34.08 ;
    RECT 75.315 33.32 75.535 34.08 ;
    RECT 76.015 33.32 76.225 34.08 ;
    RECT 76.705 33.32 76.92 34.08 ;
    RECT 77.4 33.32 77.62 34.08 ;
    RECT 78.1 33.32 78.32 34.08 ;
    RECT 78.8 33.32 79.02 34.08 ;
    RECT 79.5 33.32 81.115 34.08 ;
    RECT 81.595 33.32 81.815 34.08 ;
    RECT 82.295 33.32 82.515 34.08 ;
    RECT 82.995 33.32 83.055 34.08 ;
    RECT 83.055 33.23 83.335 34.17 ;
    RECT 83.335 33.32 83.505 34.08 ;
    RECT 26.71 32.56 26.88 33.32 ;
    RECT 26.88 32.47 27.16 33.41 ;
    RECT 27.16 32.56 27.32 33.32 ;
    RECT 27.8 32.56 28.02 33.32 ;
    RECT 28.5 32.56 28.72 33.32 ;
    RECT 29.2 32.56 30.815 33.32 ;
    RECT 31.295 32.56 31.515 33.32 ;
    RECT 31.995 32.56 32.21 33.32 ;
    RECT 32.69 32.56 32.91 33.32 ;
    RECT 33.39 32.56 33.61 33.32 ;
    RECT 34.09 32.56 34.31 33.32 ;
    RECT 34.79 32.56 35.005 33.32 ;
    RECT 35.485 32.56 36.405 33.32 ;
    RECT 36.885 32.56 37.105 33.32 ;
    RECT 37.585 32.56 37.8 33.32 ;
    RECT 38.28 32.56 38.5 33.32 ;
    RECT 38.98 32.56 39.2 33.32 ;
    RECT 39.68 32.56 39.895 33.32 ;
    RECT 40.375 32.56 40.595 33.32 ;
    RECT 41.075 32.56 41.995 33.32 ;
    RECT 42.475 32.56 42.69 33.32 ;
    RECT 43.17 32.56 43.39 33.32 ;
    RECT 43.87 32.56 44.09 33.32 ;
    RECT 44.57 32.56 44.79 33.32 ;
    RECT 45.27 32.56 45.485 33.32 ;
    RECT 45.965 32.56 46.185 33.32 ;
    RECT 46.665 32.56 47.58 33.32 ;
    RECT 48.06 32.56 48.28 33.32 ;
    RECT 48.76 32.56 48.98 33.32 ;
    RECT 49.46 32.56 49.68 33.32 ;
    RECT 50.16 32.56 50.375 33.32 ;
    RECT 50.855 32.56 51.775 33.32 ;
    RECT 52.255 32.56 53.17 33.32 ;
    RECT 53.65 32.56 53.87 33.32 ;
    RECT 54.35 32.56 54.57 33.32 ;
    RECT 55.05 32.56 55.265 33.32 ;
    RECT 55.745 32.56 55.965 33.32 ;
    RECT 56.445 32.56 56.665 33.32 ;
    RECT 57.145 32.56 58.06 33.32 ;
    RECT 58.54 32.56 59.46 33.32 ;
    RECT 59.94 32.56 60.16 33.32 ;
    RECT 60.64 32.56 60.855 33.32 ;
    RECT 61.335 32.56 61.555 33.32 ;
    RECT 62.035 32.56 62.25 33.32 ;
    RECT 62.73 32.56 63.65 33.32 ;
    RECT 64.13 32.56 64.345 33.32 ;
    RECT 64.825 32.56 65.045 33.32 ;
    RECT 65.525 32.56 65.745 33.32 ;
    RECT 66.225 32.56 66.445 33.32 ;
    RECT 66.925 32.56 67.14 33.32 ;
    RECT 67.62 32.56 67.84 33.32 ;
    RECT 68.32 32.56 69.235 33.32 ;
    RECT 69.715 32.56 69.935 33.32 ;
    RECT 70.415 32.56 70.635 33.32 ;
    RECT 71.115 32.56 71.335 33.32 ;
    RECT 71.815 32.56 72.035 33.32 ;
    RECT 72.515 32.56 72.735 33.32 ;
    RECT 73.215 32.56 73.435 33.32 ;
    RECT 73.915 32.56 74.835 33.32 ;
    RECT 75.315 32.56 75.535 33.32 ;
    RECT 76.015 32.56 76.225 33.32 ;
    RECT 76.705 32.56 76.92 33.32 ;
    RECT 77.4 32.56 77.62 33.32 ;
    RECT 78.1 32.56 78.32 33.32 ;
    RECT 78.8 32.56 79.02 33.32 ;
    RECT 79.5 32.56 81.115 33.32 ;
    RECT 81.595 32.56 81.815 33.32 ;
    RECT 82.295 32.56 82.515 33.32 ;
    RECT 82.995 32.56 83.055 33.32 ;
    RECT 83.055 32.47 83.335 33.41 ;
    RECT 83.335 32.56 83.505 33.32 ;
    RECT 26.71 31.8 26.88 32.56 ;
    RECT 26.88 31.71 27.16 32.65 ;
    RECT 27.16 31.8 27.32 32.56 ;
    RECT 27.8 31.8 28.02 32.56 ;
    RECT 28.5 31.8 28.72 32.56 ;
    RECT 29.2 31.8 30.815 32.56 ;
    RECT 31.295 31.8 31.515 32.56 ;
    RECT 31.995 31.8 32.21 32.56 ;
    RECT 32.69 31.8 32.91 32.56 ;
    RECT 33.39 31.8 33.61 32.56 ;
    RECT 34.09 31.8 34.31 32.56 ;
    RECT 34.79 31.8 35.005 32.56 ;
    RECT 35.485 31.8 36.405 32.56 ;
    RECT 36.885 31.8 37.105 32.56 ;
    RECT 37.585 31.8 37.8 32.56 ;
    RECT 38.28 31.8 38.5 32.56 ;
    RECT 38.98 31.8 39.2 32.56 ;
    RECT 39.68 31.8 39.895 32.56 ;
    RECT 40.375 31.8 40.595 32.56 ;
    RECT 41.075 31.8 41.995 32.56 ;
    RECT 42.475 31.8 42.69 32.56 ;
    RECT 43.17 31.8 43.39 32.56 ;
    RECT 43.87 31.8 44.09 32.56 ;
    RECT 44.57 31.8 44.79 32.56 ;
    RECT 45.27 31.8 45.485 32.56 ;
    RECT 45.965 31.8 46.185 32.56 ;
    RECT 46.665 31.8 47.58 32.56 ;
    RECT 48.06 31.8 48.28 32.56 ;
    RECT 48.76 31.8 48.98 32.56 ;
    RECT 49.46 31.8 49.68 32.56 ;
    RECT 50.16 31.8 50.375 32.56 ;
    RECT 50.855 31.8 51.775 32.56 ;
    RECT 52.255 31.8 53.17 32.56 ;
    RECT 53.65 31.8 53.87 32.56 ;
    RECT 54.35 31.8 54.57 32.56 ;
    RECT 55.05 31.8 55.265 32.56 ;
    RECT 55.745 31.8 55.965 32.56 ;
    RECT 56.445 31.8 56.665 32.56 ;
    RECT 57.145 31.8 58.06 32.56 ;
    RECT 58.54 31.8 59.46 32.56 ;
    RECT 59.94 31.8 60.16 32.56 ;
    RECT 60.64 31.8 60.855 32.56 ;
    RECT 61.335 31.8 61.555 32.56 ;
    RECT 62.035 31.8 62.25 32.56 ;
    RECT 62.73 31.8 63.65 32.56 ;
    RECT 64.13 31.8 64.345 32.56 ;
    RECT 64.825 31.8 65.045 32.56 ;
    RECT 65.525 31.8 65.745 32.56 ;
    RECT 66.225 31.8 66.445 32.56 ;
    RECT 66.925 31.8 67.14 32.56 ;
    RECT 67.62 31.8 67.84 32.56 ;
    RECT 68.32 31.8 69.235 32.56 ;
    RECT 69.715 31.8 69.935 32.56 ;
    RECT 70.415 31.8 70.635 32.56 ;
    RECT 71.115 31.8 71.335 32.56 ;
    RECT 71.815 31.8 72.035 32.56 ;
    RECT 72.515 31.8 72.735 32.56 ;
    RECT 73.215 31.8 73.435 32.56 ;
    RECT 73.915 31.8 74.835 32.56 ;
    RECT 75.315 31.8 75.535 32.56 ;
    RECT 76.015 31.8 76.225 32.56 ;
    RECT 76.705 31.8 76.92 32.56 ;
    RECT 77.4 31.8 77.62 32.56 ;
    RECT 78.1 31.8 78.32 32.56 ;
    RECT 78.8 31.8 79.02 32.56 ;
    RECT 79.5 31.8 81.115 32.56 ;
    RECT 81.595 31.8 81.815 32.56 ;
    RECT 82.295 31.8 82.515 32.56 ;
    RECT 82.995 31.8 83.055 32.56 ;
    RECT 83.055 31.71 83.335 32.65 ;
    RECT 83.335 31.8 83.505 32.56 ;
    RECT 26.71 31.04 26.88 31.8 ;
    RECT 26.88 30.95 27.16 31.89 ;
    RECT 27.16 31.04 27.32 31.8 ;
    RECT 27.8 31.04 28.02 31.8 ;
    RECT 28.5 31.04 28.72 31.8 ;
    RECT 29.2 31.04 30.815 31.8 ;
    RECT 31.295 31.04 31.515 31.8 ;
    RECT 31.995 31.04 32.21 31.8 ;
    RECT 32.69 31.04 32.91 31.8 ;
    RECT 33.39 31.04 33.61 31.8 ;
    RECT 34.09 31.04 34.31 31.8 ;
    RECT 34.79 31.04 35.005 31.8 ;
    RECT 35.485 31.04 36.405 31.8 ;
    RECT 36.885 31.04 37.105 31.8 ;
    RECT 37.585 31.04 37.8 31.8 ;
    RECT 38.28 31.04 38.5 31.8 ;
    RECT 38.98 31.04 39.2 31.8 ;
    RECT 39.68 31.04 39.895 31.8 ;
    RECT 40.375 31.04 40.595 31.8 ;
    RECT 41.075 31.04 41.995 31.8 ;
    RECT 42.475 31.04 42.69 31.8 ;
    RECT 43.17 31.04 43.39 31.8 ;
    RECT 43.87 31.04 44.09 31.8 ;
    RECT 44.57 31.04 44.79 31.8 ;
    RECT 45.27 31.04 45.485 31.8 ;
    RECT 45.965 31.04 46.185 31.8 ;
    RECT 46.665 31.04 47.58 31.8 ;
    RECT 48.06 31.04 48.28 31.8 ;
    RECT 48.76 31.04 48.98 31.8 ;
    RECT 49.46 31.04 49.68 31.8 ;
    RECT 50.16 31.04 50.375 31.8 ;
    RECT 50.855 31.04 51.775 31.8 ;
    RECT 52.255 31.04 53.17 31.8 ;
    RECT 53.65 31.04 53.87 31.8 ;
    RECT 54.35 31.04 54.57 31.8 ;
    RECT 55.05 31.04 55.265 31.8 ;
    RECT 55.745 31.04 55.965 31.8 ;
    RECT 56.445 31.04 56.665 31.8 ;
    RECT 57.145 31.04 58.06 31.8 ;
    RECT 58.54 31.04 59.46 31.8 ;
    RECT 59.94 31.04 60.16 31.8 ;
    RECT 60.64 31.04 60.855 31.8 ;
    RECT 61.335 31.04 61.555 31.8 ;
    RECT 62.035 31.04 62.25 31.8 ;
    RECT 62.73 31.04 63.65 31.8 ;
    RECT 64.13 31.04 64.345 31.8 ;
    RECT 64.825 31.04 65.045 31.8 ;
    RECT 65.525 31.04 65.745 31.8 ;
    RECT 66.225 31.04 66.445 31.8 ;
    RECT 66.925 31.04 67.14 31.8 ;
    RECT 67.62 31.04 67.84 31.8 ;
    RECT 68.32 31.04 69.235 31.8 ;
    RECT 69.715 31.04 69.935 31.8 ;
    RECT 70.415 31.04 70.635 31.8 ;
    RECT 71.115 31.04 71.335 31.8 ;
    RECT 71.815 31.04 72.035 31.8 ;
    RECT 72.515 31.04 72.735 31.8 ;
    RECT 73.215 31.04 73.435 31.8 ;
    RECT 73.915 31.04 74.835 31.8 ;
    RECT 75.315 31.04 75.535 31.8 ;
    RECT 76.015 31.04 76.225 31.8 ;
    RECT 76.705 31.04 76.92 31.8 ;
    RECT 77.4 31.04 77.62 31.8 ;
    RECT 78.1 31.04 78.32 31.8 ;
    RECT 78.8 31.04 79.02 31.8 ;
    RECT 79.5 31.04 81.115 31.8 ;
    RECT 81.595 31.04 81.815 31.8 ;
    RECT 82.295 31.04 82.515 31.8 ;
    RECT 82.995 31.04 83.055 31.8 ;
    RECT 83.055 30.95 83.335 31.89 ;
    RECT 83.335 31.04 83.505 31.8 ;
    RECT 26.71 30.28 26.88 31.04 ;
    RECT 26.88 30.19 27.16 31.13 ;
    RECT 27.16 30.28 27.32 31.04 ;
    RECT 27.8 30.28 28.02 31.04 ;
    RECT 28.5 30.28 28.72 31.04 ;
    RECT 29.2 30.28 30.815 31.04 ;
    RECT 31.295 30.28 31.515 31.04 ;
    RECT 31.995 30.28 32.21 31.04 ;
    RECT 32.69 30.28 32.91 31.04 ;
    RECT 33.39 30.28 33.61 31.04 ;
    RECT 34.09 30.28 34.31 31.04 ;
    RECT 34.79 30.28 35.005 31.04 ;
    RECT 35.485 30.28 36.405 31.04 ;
    RECT 36.885 30.28 37.105 31.04 ;
    RECT 37.585 30.28 37.8 31.04 ;
    RECT 38.28 30.28 38.5 31.04 ;
    RECT 38.98 30.28 39.2 31.04 ;
    RECT 39.68 30.28 39.895 31.04 ;
    RECT 40.375 30.28 40.595 31.04 ;
    RECT 41.075 30.28 41.995 31.04 ;
    RECT 42.475 30.28 42.69 31.04 ;
    RECT 43.17 30.28 43.39 31.04 ;
    RECT 43.87 30.28 44.09 31.04 ;
    RECT 44.57 30.28 44.79 31.04 ;
    RECT 45.27 30.28 45.485 31.04 ;
    RECT 45.965 30.28 46.185 31.04 ;
    RECT 46.665 30.28 47.58 31.04 ;
    RECT 48.06 30.28 48.28 31.04 ;
    RECT 48.76 30.28 48.98 31.04 ;
    RECT 49.46 30.28 49.68 31.04 ;
    RECT 50.16 30.28 50.375 31.04 ;
    RECT 50.855 30.28 51.775 31.04 ;
    RECT 52.255 30.28 53.17 31.04 ;
    RECT 53.65 30.28 53.87 31.04 ;
    RECT 54.35 30.28 54.57 31.04 ;
    RECT 55.05 30.28 55.265 31.04 ;
    RECT 55.745 30.28 55.965 31.04 ;
    RECT 56.445 30.28 56.665 31.04 ;
    RECT 57.145 30.28 58.06 31.04 ;
    RECT 58.54 30.28 59.46 31.04 ;
    RECT 59.94 30.28 60.16 31.04 ;
    RECT 60.64 30.28 60.855 31.04 ;
    RECT 61.335 30.28 61.555 31.04 ;
    RECT 62.035 30.28 62.25 31.04 ;
    RECT 62.73 30.28 63.65 31.04 ;
    RECT 64.13 30.28 64.345 31.04 ;
    RECT 64.825 30.28 65.045 31.04 ;
    RECT 65.525 30.28 65.745 31.04 ;
    RECT 66.225 30.28 66.445 31.04 ;
    RECT 66.925 30.28 67.14 31.04 ;
    RECT 67.62 30.28 67.84 31.04 ;
    RECT 68.32 30.28 69.235 31.04 ;
    RECT 69.715 30.28 69.935 31.04 ;
    RECT 70.415 30.28 70.635 31.04 ;
    RECT 71.115 30.28 71.335 31.04 ;
    RECT 71.815 30.28 72.035 31.04 ;
    RECT 72.515 30.28 72.735 31.04 ;
    RECT 73.215 30.28 73.435 31.04 ;
    RECT 73.915 30.28 74.835 31.04 ;
    RECT 75.315 30.28 75.535 31.04 ;
    RECT 76.015 30.28 76.225 31.04 ;
    RECT 76.705 30.28 76.92 31.04 ;
    RECT 77.4 30.28 77.62 31.04 ;
    RECT 78.1 30.28 78.32 31.04 ;
    RECT 78.8 30.28 79.02 31.04 ;
    RECT 79.5 30.28 81.115 31.04 ;
    RECT 81.595 30.28 81.815 31.04 ;
    RECT 82.295 30.28 82.515 31.04 ;
    RECT 82.995 30.28 83.055 31.04 ;
    RECT 83.055 30.19 83.335 31.13 ;
    RECT 83.335 30.28 83.505 31.04 ;
    RECT 26.71 29.52 26.88 30.28 ;
    RECT 26.88 29.43 27.16 30.37 ;
    RECT 27.16 29.52 27.32 30.28 ;
    RECT 27.8 29.52 28.02 30.28 ;
    RECT 28.5 29.52 28.72 30.28 ;
    RECT 29.2 29.52 30.815 30.28 ;
    RECT 31.295 29.52 31.515 30.28 ;
    RECT 31.995 29.52 32.21 30.28 ;
    RECT 32.69 29.52 32.91 30.28 ;
    RECT 33.39 29.52 33.61 30.28 ;
    RECT 34.09 29.52 34.31 30.28 ;
    RECT 34.79 29.52 35.005 30.28 ;
    RECT 35.485 29.52 36.405 30.28 ;
    RECT 36.885 29.52 37.105 30.28 ;
    RECT 37.585 29.52 37.8 30.28 ;
    RECT 38.28 29.52 38.5 30.28 ;
    RECT 38.98 29.52 39.2 30.28 ;
    RECT 39.68 29.52 39.895 30.28 ;
    RECT 40.375 29.52 40.595 30.28 ;
    RECT 41.075 29.52 41.995 30.28 ;
    RECT 42.475 29.52 42.69 30.28 ;
    RECT 43.17 29.52 43.39 30.28 ;
    RECT 43.87 29.52 44.09 30.28 ;
    RECT 44.57 29.52 44.79 30.28 ;
    RECT 45.27 29.52 45.485 30.28 ;
    RECT 45.965 29.52 46.185 30.28 ;
    RECT 46.665 29.52 47.58 30.28 ;
    RECT 48.06 29.52 48.28 30.28 ;
    RECT 48.76 29.52 48.98 30.28 ;
    RECT 49.46 29.52 49.68 30.28 ;
    RECT 50.16 29.52 50.375 30.28 ;
    RECT 50.855 29.52 51.775 30.28 ;
    RECT 52.255 29.52 53.17 30.28 ;
    RECT 53.65 29.52 53.87 30.28 ;
    RECT 54.35 29.52 54.57 30.28 ;
    RECT 55.05 29.52 55.265 30.28 ;
    RECT 55.745 29.52 55.965 30.28 ;
    RECT 56.445 29.52 56.665 30.28 ;
    RECT 57.145 29.52 58.06 30.28 ;
    RECT 58.54 29.52 59.46 30.28 ;
    RECT 59.94 29.52 60.16 30.28 ;
    RECT 60.64 29.52 60.855 30.28 ;
    RECT 61.335 29.52 61.555 30.28 ;
    RECT 62.035 29.52 62.25 30.28 ;
    RECT 62.73 29.52 63.65 30.28 ;
    RECT 64.13 29.52 64.345 30.28 ;
    RECT 64.825 29.52 65.045 30.28 ;
    RECT 65.525 29.52 65.745 30.28 ;
    RECT 66.225 29.52 66.445 30.28 ;
    RECT 66.925 29.52 67.14 30.28 ;
    RECT 67.62 29.52 67.84 30.28 ;
    RECT 68.32 29.52 69.235 30.28 ;
    RECT 69.715 29.52 69.935 30.28 ;
    RECT 70.415 29.52 70.635 30.28 ;
    RECT 71.115 29.52 71.335 30.28 ;
    RECT 71.815 29.52 72.035 30.28 ;
    RECT 72.515 29.52 72.735 30.28 ;
    RECT 73.215 29.52 73.435 30.28 ;
    RECT 73.915 29.52 74.835 30.28 ;
    RECT 75.315 29.52 75.535 30.28 ;
    RECT 76.015 29.52 76.225 30.28 ;
    RECT 76.705 29.52 76.92 30.28 ;
    RECT 77.4 29.52 77.62 30.28 ;
    RECT 78.1 29.52 78.32 30.28 ;
    RECT 78.8 29.52 79.02 30.28 ;
    RECT 79.5 29.52 81.115 30.28 ;
    RECT 81.595 29.52 81.815 30.28 ;
    RECT 82.295 29.52 82.515 30.28 ;
    RECT 82.995 29.52 83.055 30.28 ;
    RECT 83.055 29.43 83.335 30.37 ;
    RECT 83.335 29.52 83.505 30.28 ;
    RECT 26.71 28.76 26.88 29.52 ;
    RECT 26.88 28.67 27.16 29.61 ;
    RECT 27.16 28.76 27.32 29.52 ;
    RECT 27.8 28.76 28.02 29.52 ;
    RECT 28.5 28.76 28.72 29.52 ;
    RECT 29.2 28.76 30.815 29.52 ;
    RECT 31.295 28.76 31.515 29.52 ;
    RECT 31.995 28.76 32.21 29.52 ;
    RECT 32.69 28.76 32.91 29.52 ;
    RECT 33.39 28.76 33.61 29.52 ;
    RECT 34.09 28.76 34.31 29.52 ;
    RECT 34.79 28.76 35.005 29.52 ;
    RECT 35.485 28.76 36.405 29.52 ;
    RECT 36.885 28.76 37.105 29.52 ;
    RECT 37.585 28.76 37.8 29.52 ;
    RECT 38.28 28.76 38.5 29.52 ;
    RECT 38.98 28.76 39.2 29.52 ;
    RECT 39.68 28.76 39.895 29.52 ;
    RECT 40.375 28.76 40.595 29.52 ;
    RECT 41.075 28.76 41.995 29.52 ;
    RECT 42.475 28.76 42.69 29.52 ;
    RECT 43.17 28.76 43.39 29.52 ;
    RECT 43.87 28.76 44.09 29.52 ;
    RECT 44.57 28.76 44.79 29.52 ;
    RECT 45.27 28.76 45.485 29.52 ;
    RECT 45.965 28.76 46.185 29.52 ;
    RECT 46.665 28.76 47.58 29.52 ;
    RECT 48.06 28.76 48.28 29.52 ;
    RECT 48.76 28.76 48.98 29.52 ;
    RECT 49.46 28.76 49.68 29.52 ;
    RECT 50.16 28.76 50.375 29.52 ;
    RECT 50.855 28.76 51.775 29.52 ;
    RECT 52.255 28.76 53.17 29.52 ;
    RECT 53.65 28.76 53.87 29.52 ;
    RECT 54.35 28.76 54.57 29.52 ;
    RECT 55.05 28.76 55.265 29.52 ;
    RECT 55.745 28.76 55.965 29.52 ;
    RECT 56.445 28.76 56.665 29.52 ;
    RECT 57.145 28.76 58.06 29.52 ;
    RECT 58.54 28.76 59.46 29.52 ;
    RECT 59.94 28.76 60.16 29.52 ;
    RECT 60.64 28.76 60.855 29.52 ;
    RECT 61.335 28.76 61.555 29.52 ;
    RECT 62.035 28.76 62.25 29.52 ;
    RECT 62.73 28.76 63.65 29.52 ;
    RECT 64.13 28.76 64.345 29.52 ;
    RECT 64.825 28.76 65.045 29.52 ;
    RECT 65.525 28.76 65.745 29.52 ;
    RECT 66.225 28.76 66.445 29.52 ;
    RECT 66.925 28.76 67.14 29.52 ;
    RECT 67.62 28.76 67.84 29.52 ;
    RECT 68.32 28.76 69.235 29.52 ;
    RECT 69.715 28.76 69.935 29.52 ;
    RECT 70.415 28.76 70.635 29.52 ;
    RECT 71.115 28.76 71.335 29.52 ;
    RECT 71.815 28.76 72.035 29.52 ;
    RECT 72.515 28.76 72.735 29.52 ;
    RECT 73.215 28.76 73.435 29.52 ;
    RECT 73.915 28.76 74.835 29.52 ;
    RECT 75.315 28.76 75.535 29.52 ;
    RECT 76.015 28.76 76.225 29.52 ;
    RECT 76.705 28.76 76.92 29.52 ;
    RECT 77.4 28.76 77.62 29.52 ;
    RECT 78.1 28.76 78.32 29.52 ;
    RECT 78.8 28.76 79.02 29.52 ;
    RECT 79.5 28.76 81.115 29.52 ;
    RECT 81.595 28.76 81.815 29.52 ;
    RECT 82.295 28.76 82.515 29.52 ;
    RECT 82.995 28.76 83.055 29.52 ;
    RECT 83.055 28.67 83.335 29.61 ;
    RECT 83.335 28.76 83.505 29.52 ;
    RECT 26.71 28.0 26.88 28.76 ;
    RECT 26.88 27.91 27.16 28.85 ;
    RECT 27.16 28.0 27.32 28.76 ;
    RECT 27.8 28.0 28.02 28.76 ;
    RECT 28.5 28.0 28.72 28.76 ;
    RECT 29.2 28.0 30.815 28.76 ;
    RECT 31.295 28.0 31.515 28.76 ;
    RECT 31.995 28.0 32.21 28.76 ;
    RECT 32.69 28.0 32.91 28.76 ;
    RECT 33.39 28.0 33.61 28.76 ;
    RECT 34.09 28.0 34.31 28.76 ;
    RECT 34.79 28.0 35.005 28.76 ;
    RECT 35.485 28.0 36.405 28.76 ;
    RECT 36.885 28.0 37.105 28.76 ;
    RECT 37.585 28.0 37.8 28.76 ;
    RECT 38.28 28.0 38.5 28.76 ;
    RECT 38.98 28.0 39.2 28.76 ;
    RECT 39.68 28.0 39.895 28.76 ;
    RECT 40.375 28.0 40.595 28.76 ;
    RECT 41.075 28.0 41.995 28.76 ;
    RECT 42.475 28.0 42.69 28.76 ;
    RECT 43.17 28.0 43.39 28.76 ;
    RECT 43.87 28.0 44.09 28.76 ;
    RECT 44.57 28.0 44.79 28.76 ;
    RECT 45.27 28.0 45.485 28.76 ;
    RECT 45.965 28.0 46.185 28.76 ;
    RECT 46.665 28.0 47.58 28.76 ;
    RECT 48.06 28.0 48.28 28.76 ;
    RECT 48.76 28.0 48.98 28.76 ;
    RECT 49.46 28.0 49.68 28.76 ;
    RECT 50.16 28.0 50.375 28.76 ;
    RECT 50.855 28.0 51.775 28.76 ;
    RECT 52.255 28.0 53.17 28.76 ;
    RECT 53.65 28.0 53.87 28.76 ;
    RECT 54.35 28.0 54.57 28.76 ;
    RECT 55.05 28.0 55.265 28.76 ;
    RECT 55.745 28.0 55.965 28.76 ;
    RECT 56.445 28.0 56.665 28.76 ;
    RECT 57.145 28.0 58.06 28.76 ;
    RECT 58.54 28.0 59.46 28.76 ;
    RECT 59.94 28.0 60.16 28.76 ;
    RECT 60.64 28.0 60.855 28.76 ;
    RECT 61.335 28.0 61.555 28.76 ;
    RECT 62.035 28.0 62.25 28.76 ;
    RECT 62.73 28.0 63.65 28.76 ;
    RECT 64.13 28.0 64.345 28.76 ;
    RECT 64.825 28.0 65.045 28.76 ;
    RECT 65.525 28.0 65.745 28.76 ;
    RECT 66.225 28.0 66.445 28.76 ;
    RECT 66.925 28.0 67.14 28.76 ;
    RECT 67.62 28.0 67.84 28.76 ;
    RECT 68.32 28.0 69.235 28.76 ;
    RECT 69.715 28.0 69.935 28.76 ;
    RECT 70.415 28.0 70.635 28.76 ;
    RECT 71.115 28.0 71.335 28.76 ;
    RECT 71.815 28.0 72.035 28.76 ;
    RECT 72.515 28.0 72.735 28.76 ;
    RECT 73.215 28.0 73.435 28.76 ;
    RECT 73.915 28.0 74.835 28.76 ;
    RECT 75.315 28.0 75.535 28.76 ;
    RECT 76.015 28.0 76.225 28.76 ;
    RECT 76.705 28.0 76.92 28.76 ;
    RECT 77.4 28.0 77.62 28.76 ;
    RECT 78.1 28.0 78.32 28.76 ;
    RECT 78.8 28.0 79.02 28.76 ;
    RECT 79.5 28.0 81.115 28.76 ;
    RECT 81.595 28.0 81.815 28.76 ;
    RECT 82.295 28.0 82.515 28.76 ;
    RECT 82.995 28.0 83.055 28.76 ;
    RECT 83.055 27.91 83.335 28.85 ;
    RECT 83.335 28.0 83.505 28.76 ;
    RECT 26.71 27.24 26.88 28.0 ;
    RECT 26.88 27.15 27.16 28.09 ;
    RECT 27.16 27.24 27.32 28.0 ;
    RECT 27.8 27.24 28.02 28.0 ;
    RECT 28.5 27.24 28.72 28.0 ;
    RECT 29.2 27.24 30.815 28.0 ;
    RECT 31.295 27.24 31.515 28.0 ;
    RECT 31.995 27.24 32.21 28.0 ;
    RECT 32.69 27.24 32.91 28.0 ;
    RECT 33.39 27.24 33.61 28.0 ;
    RECT 34.09 27.24 34.31 28.0 ;
    RECT 34.79 27.24 35.005 28.0 ;
    RECT 35.485 27.24 36.405 28.0 ;
    RECT 36.885 27.24 37.105 28.0 ;
    RECT 37.585 27.24 37.8 28.0 ;
    RECT 38.28 27.24 38.5 28.0 ;
    RECT 38.98 27.24 39.2 28.0 ;
    RECT 39.68 27.24 39.895 28.0 ;
    RECT 40.375 27.24 40.595 28.0 ;
    RECT 41.075 27.24 41.995 28.0 ;
    RECT 42.475 27.24 42.69 28.0 ;
    RECT 43.17 27.24 43.39 28.0 ;
    RECT 43.87 27.24 44.09 28.0 ;
    RECT 44.57 27.24 44.79 28.0 ;
    RECT 45.27 27.24 45.485 28.0 ;
    RECT 45.965 27.24 46.185 28.0 ;
    RECT 46.665 27.24 47.58 28.0 ;
    RECT 48.06 27.24 48.28 28.0 ;
    RECT 48.76 27.24 48.98 28.0 ;
    RECT 49.46 27.24 49.68 28.0 ;
    RECT 50.16 27.24 50.375 28.0 ;
    RECT 50.855 27.24 51.775 28.0 ;
    RECT 52.255 27.24 53.17 28.0 ;
    RECT 53.65 27.24 53.87 28.0 ;
    RECT 54.35 27.24 54.57 28.0 ;
    RECT 55.05 27.24 55.265 28.0 ;
    RECT 55.745 27.24 55.965 28.0 ;
    RECT 56.445 27.24 56.665 28.0 ;
    RECT 57.145 27.24 58.06 28.0 ;
    RECT 58.54 27.24 59.46 28.0 ;
    RECT 59.94 27.24 60.16 28.0 ;
    RECT 60.64 27.24 60.855 28.0 ;
    RECT 61.335 27.24 61.555 28.0 ;
    RECT 62.035 27.24 62.25 28.0 ;
    RECT 62.73 27.24 63.65 28.0 ;
    RECT 64.13 27.24 64.345 28.0 ;
    RECT 64.825 27.24 65.045 28.0 ;
    RECT 65.525 27.24 65.745 28.0 ;
    RECT 66.225 27.24 66.445 28.0 ;
    RECT 66.925 27.24 67.14 28.0 ;
    RECT 67.62 27.24 67.84 28.0 ;
    RECT 68.32 27.24 69.235 28.0 ;
    RECT 69.715 27.24 69.935 28.0 ;
    RECT 70.415 27.24 70.635 28.0 ;
    RECT 71.115 27.24 71.335 28.0 ;
    RECT 71.815 27.24 72.035 28.0 ;
    RECT 72.515 27.24 72.735 28.0 ;
    RECT 73.215 27.24 73.435 28.0 ;
    RECT 73.915 27.24 74.835 28.0 ;
    RECT 75.315 27.24 75.535 28.0 ;
    RECT 76.015 27.24 76.225 28.0 ;
    RECT 76.705 27.24 76.92 28.0 ;
    RECT 77.4 27.24 77.62 28.0 ;
    RECT 78.1 27.24 78.32 28.0 ;
    RECT 78.8 27.24 79.02 28.0 ;
    RECT 79.5 27.24 81.115 28.0 ;
    RECT 81.595 27.24 81.815 28.0 ;
    RECT 82.295 27.24 82.515 28.0 ;
    RECT 82.995 27.24 83.055 28.0 ;
    RECT 83.055 27.15 83.335 28.09 ;
    RECT 83.335 27.24 83.505 28.0 ;
    RECT 26.71 26.48 26.88 27.24 ;
    RECT 26.88 26.39 27.16 27.33 ;
    RECT 27.16 26.48 27.32 27.24 ;
    RECT 27.8 26.48 28.02 27.24 ;
    RECT 28.5 26.48 28.72 27.24 ;
    RECT 29.2 26.48 30.815 27.24 ;
    RECT 31.295 26.48 31.515 27.24 ;
    RECT 31.995 26.48 32.21 27.24 ;
    RECT 32.69 26.48 32.91 27.24 ;
    RECT 33.39 26.48 33.61 27.24 ;
    RECT 34.09 26.48 34.31 27.24 ;
    RECT 34.79 26.48 35.005 27.24 ;
    RECT 35.485 26.48 36.405 27.24 ;
    RECT 36.885 26.48 37.105 27.24 ;
    RECT 37.585 26.48 37.8 27.24 ;
    RECT 38.28 26.48 38.5 27.24 ;
    RECT 38.98 26.48 39.2 27.24 ;
    RECT 39.68 26.48 39.895 27.24 ;
    RECT 40.375 26.48 40.595 27.24 ;
    RECT 41.075 26.48 41.995 27.24 ;
    RECT 42.475 26.48 42.69 27.24 ;
    RECT 43.17 26.48 43.39 27.24 ;
    RECT 43.87 26.48 44.09 27.24 ;
    RECT 44.57 26.48 44.79 27.24 ;
    RECT 45.27 26.48 45.485 27.24 ;
    RECT 45.965 26.48 46.185 27.24 ;
    RECT 46.665 26.48 47.58 27.24 ;
    RECT 48.06 26.48 48.28 27.24 ;
    RECT 48.76 26.48 48.98 27.24 ;
    RECT 49.46 26.48 49.68 27.24 ;
    RECT 50.16 26.48 50.375 27.24 ;
    RECT 50.855 26.48 51.775 27.24 ;
    RECT 52.255 26.48 53.17 27.24 ;
    RECT 53.65 26.48 53.87 27.24 ;
    RECT 54.35 26.48 54.57 27.24 ;
    RECT 55.05 26.48 55.265 27.24 ;
    RECT 55.745 26.48 55.965 27.24 ;
    RECT 56.445 26.48 56.665 27.24 ;
    RECT 57.145 26.48 58.06 27.24 ;
    RECT 58.54 26.48 59.46 27.24 ;
    RECT 59.94 26.48 60.16 27.24 ;
    RECT 60.64 26.48 60.855 27.24 ;
    RECT 61.335 26.48 61.555 27.24 ;
    RECT 62.035 26.48 62.25 27.24 ;
    RECT 62.73 26.48 63.65 27.24 ;
    RECT 64.13 26.48 64.345 27.24 ;
    RECT 64.825 26.48 65.045 27.24 ;
    RECT 65.525 26.48 65.745 27.24 ;
    RECT 66.225 26.48 66.445 27.24 ;
    RECT 66.925 26.48 67.14 27.24 ;
    RECT 67.62 26.48 67.84 27.24 ;
    RECT 68.32 26.48 69.235 27.24 ;
    RECT 69.715 26.48 69.935 27.24 ;
    RECT 70.415 26.48 70.635 27.24 ;
    RECT 71.115 26.48 71.335 27.24 ;
    RECT 71.815 26.48 72.035 27.24 ;
    RECT 72.515 26.48 72.735 27.24 ;
    RECT 73.215 26.48 73.435 27.24 ;
    RECT 73.915 26.48 74.835 27.24 ;
    RECT 75.315 26.48 75.535 27.24 ;
    RECT 76.015 26.48 76.225 27.24 ;
    RECT 76.705 26.48 76.92 27.24 ;
    RECT 77.4 26.48 77.62 27.24 ;
    RECT 78.1 26.48 78.32 27.24 ;
    RECT 78.8 26.48 79.02 27.24 ;
    RECT 79.5 26.48 81.115 27.24 ;
    RECT 81.595 26.48 81.815 27.24 ;
    RECT 82.295 26.48 82.515 27.24 ;
    RECT 82.995 26.48 83.055 27.24 ;
    RECT 83.055 26.39 83.335 27.33 ;
    RECT 83.335 26.48 83.505 27.24 ;
    RECT 26.71 25.72 26.88 26.48 ;
    RECT 26.88 25.63 27.16 26.57 ;
    RECT 27.16 25.72 27.32 26.48 ;
    RECT 27.8 25.72 28.02 26.48 ;
    RECT 28.5 25.72 28.72 26.48 ;
    RECT 29.2 25.72 30.815 26.48 ;
    RECT 31.295 25.72 31.515 26.48 ;
    RECT 31.995 25.72 32.21 26.48 ;
    RECT 32.69 25.72 32.91 26.48 ;
    RECT 33.39 25.72 33.61 26.48 ;
    RECT 34.09 25.72 34.31 26.48 ;
    RECT 34.79 25.72 35.005 26.48 ;
    RECT 35.485 25.72 36.405 26.48 ;
    RECT 36.885 25.72 37.105 26.48 ;
    RECT 37.585 25.72 37.8 26.48 ;
    RECT 38.28 25.72 38.5 26.48 ;
    RECT 38.98 25.72 39.2 26.48 ;
    RECT 39.68 25.72 39.895 26.48 ;
    RECT 40.375 25.72 40.595 26.48 ;
    RECT 41.075 25.72 41.995 26.48 ;
    RECT 42.475 25.72 42.69 26.48 ;
    RECT 43.17 25.72 43.39 26.48 ;
    RECT 43.87 25.72 44.09 26.48 ;
    RECT 44.57 25.72 44.79 26.48 ;
    RECT 45.27 25.72 45.485 26.48 ;
    RECT 45.965 25.72 46.185 26.48 ;
    RECT 46.665 25.72 47.58 26.48 ;
    RECT 48.06 25.72 48.28 26.48 ;
    RECT 48.76 25.72 48.98 26.48 ;
    RECT 49.46 25.72 49.68 26.48 ;
    RECT 50.16 25.72 50.375 26.48 ;
    RECT 50.855 25.72 51.775 26.48 ;
    RECT 52.255 25.72 53.17 26.48 ;
    RECT 53.65 25.72 53.87 26.48 ;
    RECT 54.35 25.72 54.57 26.48 ;
    RECT 55.05 25.72 55.265 26.48 ;
    RECT 55.745 25.72 55.965 26.48 ;
    RECT 56.445 25.72 56.665 26.48 ;
    RECT 57.145 25.72 58.06 26.48 ;
    RECT 58.54 25.72 59.46 26.48 ;
    RECT 59.94 25.72 60.16 26.48 ;
    RECT 60.64 25.72 60.855 26.48 ;
    RECT 61.335 25.72 61.555 26.48 ;
    RECT 62.035 25.72 62.25 26.48 ;
    RECT 62.73 25.72 63.65 26.48 ;
    RECT 64.13 25.72 64.345 26.48 ;
    RECT 64.825 25.72 65.045 26.48 ;
    RECT 65.525 25.72 65.745 26.48 ;
    RECT 66.225 25.72 66.445 26.48 ;
    RECT 66.925 25.72 67.14 26.48 ;
    RECT 67.62 25.72 67.84 26.48 ;
    RECT 68.32 25.72 69.235 26.48 ;
    RECT 69.715 25.72 69.935 26.48 ;
    RECT 70.415 25.72 70.635 26.48 ;
    RECT 71.115 25.72 71.335 26.48 ;
    RECT 71.815 25.72 72.035 26.48 ;
    RECT 72.515 25.72 72.735 26.48 ;
    RECT 73.215 25.72 73.435 26.48 ;
    RECT 73.915 25.72 74.835 26.48 ;
    RECT 75.315 25.72 75.535 26.48 ;
    RECT 76.015 25.72 76.225 26.48 ;
    RECT 76.705 25.72 76.92 26.48 ;
    RECT 77.4 25.72 77.62 26.48 ;
    RECT 78.1 25.72 78.32 26.48 ;
    RECT 78.8 25.72 79.02 26.48 ;
    RECT 79.5 25.72 81.115 26.48 ;
    RECT 81.595 25.72 81.815 26.48 ;
    RECT 82.295 25.72 82.515 26.48 ;
    RECT 82.995 25.72 83.055 26.48 ;
    RECT 83.055 25.63 83.335 26.57 ;
    RECT 83.335 25.72 83.505 26.48 ;
    RECT 26.71 24.96 26.88 25.72 ;
    RECT 26.88 24.87 27.16 25.81 ;
    RECT 27.16 24.96 27.32 25.72 ;
    RECT 27.8 24.96 28.02 25.72 ;
    RECT 28.5 24.96 28.72 25.72 ;
    RECT 29.2 24.96 30.815 25.72 ;
    RECT 31.295 24.96 31.515 25.72 ;
    RECT 31.995 24.96 32.21 25.72 ;
    RECT 32.69 24.96 32.91 25.72 ;
    RECT 33.39 24.96 33.61 25.72 ;
    RECT 34.09 24.96 34.31 25.72 ;
    RECT 34.79 24.96 35.005 25.72 ;
    RECT 35.485 24.96 36.405 25.72 ;
    RECT 36.885 24.96 37.105 25.72 ;
    RECT 37.585 24.96 37.8 25.72 ;
    RECT 38.28 24.96 38.5 25.72 ;
    RECT 38.98 24.96 39.2 25.72 ;
    RECT 39.68 24.96 39.895 25.72 ;
    RECT 40.375 24.96 40.595 25.72 ;
    RECT 41.075 24.96 41.995 25.72 ;
    RECT 42.475 24.96 42.69 25.72 ;
    RECT 43.17 24.96 43.39 25.72 ;
    RECT 43.87 24.96 44.09 25.72 ;
    RECT 44.57 24.96 44.79 25.72 ;
    RECT 45.27 24.96 45.485 25.72 ;
    RECT 45.965 24.96 46.185 25.72 ;
    RECT 46.665 24.96 47.58 25.72 ;
    RECT 48.06 24.96 48.28 25.72 ;
    RECT 48.76 24.96 48.98 25.72 ;
    RECT 49.46 24.96 49.68 25.72 ;
    RECT 50.16 24.96 50.375 25.72 ;
    RECT 50.855 24.96 51.775 25.72 ;
    RECT 52.255 24.96 53.17 25.72 ;
    RECT 53.65 24.96 53.87 25.72 ;
    RECT 54.35 24.96 54.57 25.72 ;
    RECT 55.05 24.96 55.265 25.72 ;
    RECT 55.745 24.96 55.965 25.72 ;
    RECT 56.445 24.96 56.665 25.72 ;
    RECT 57.145 24.96 58.06 25.72 ;
    RECT 58.54 24.96 59.46 25.72 ;
    RECT 59.94 24.96 60.16 25.72 ;
    RECT 60.64 24.96 60.855 25.72 ;
    RECT 61.335 24.96 61.555 25.72 ;
    RECT 62.035 24.96 62.25 25.72 ;
    RECT 62.73 24.96 63.65 25.72 ;
    RECT 64.13 24.96 64.345 25.72 ;
    RECT 64.825 24.96 65.045 25.72 ;
    RECT 65.525 24.96 65.745 25.72 ;
    RECT 66.225 24.96 66.445 25.72 ;
    RECT 66.925 24.96 67.14 25.72 ;
    RECT 67.62 24.96 67.84 25.72 ;
    RECT 68.32 24.96 69.235 25.72 ;
    RECT 69.715 24.96 69.935 25.72 ;
    RECT 70.415 24.96 70.635 25.72 ;
    RECT 71.115 24.96 71.335 25.72 ;
    RECT 71.815 24.96 72.035 25.72 ;
    RECT 72.515 24.96 72.735 25.72 ;
    RECT 73.215 24.96 73.435 25.72 ;
    RECT 73.915 24.96 74.835 25.72 ;
    RECT 75.315 24.96 75.535 25.72 ;
    RECT 76.015 24.96 76.225 25.72 ;
    RECT 76.705 24.96 76.92 25.72 ;
    RECT 77.4 24.96 77.62 25.72 ;
    RECT 78.1 24.96 78.32 25.72 ;
    RECT 78.8 24.96 79.02 25.72 ;
    RECT 79.5 24.96 81.115 25.72 ;
    RECT 81.595 24.96 81.815 25.72 ;
    RECT 82.295 24.96 82.515 25.72 ;
    RECT 82.995 24.96 83.055 25.72 ;
    RECT 83.055 24.87 83.335 25.81 ;
    RECT 83.335 24.96 83.505 25.72 ;
    RECT 26.71 24.2 26.88 24.96 ;
    RECT 26.88 24.11 27.16 25.05 ;
    RECT 27.16 24.2 27.32 24.96 ;
    RECT 27.8 24.2 28.02 24.96 ;
    RECT 28.5 24.2 28.72 24.96 ;
    RECT 29.2 24.2 30.815 24.96 ;
    RECT 31.295 24.2 31.515 24.96 ;
    RECT 31.995 24.2 32.21 24.96 ;
    RECT 32.69 24.2 32.91 24.96 ;
    RECT 33.39 24.2 33.61 24.96 ;
    RECT 34.09 24.2 34.31 24.96 ;
    RECT 34.79 24.2 35.005 24.96 ;
    RECT 35.485 24.2 36.405 24.96 ;
    RECT 36.885 24.2 37.105 24.96 ;
    RECT 37.585 24.2 37.8 24.96 ;
    RECT 38.28 24.2 38.5 24.96 ;
    RECT 38.98 24.2 39.2 24.96 ;
    RECT 39.68 24.2 39.895 24.96 ;
    RECT 40.375 24.2 40.595 24.96 ;
    RECT 41.075 24.2 41.995 24.96 ;
    RECT 42.475 24.2 42.69 24.96 ;
    RECT 43.17 24.2 43.39 24.96 ;
    RECT 43.87 24.2 44.09 24.96 ;
    RECT 44.57 24.2 44.79 24.96 ;
    RECT 45.27 24.2 45.485 24.96 ;
    RECT 45.965 24.2 46.185 24.96 ;
    RECT 46.665 24.2 47.58 24.96 ;
    RECT 48.06 24.2 48.28 24.96 ;
    RECT 48.76 24.2 48.98 24.96 ;
    RECT 49.46 24.2 49.68 24.96 ;
    RECT 50.16 24.2 50.375 24.96 ;
    RECT 50.855 24.2 51.775 24.96 ;
    RECT 52.255 24.2 53.17 24.96 ;
    RECT 53.65 24.2 53.87 24.96 ;
    RECT 54.35 24.2 54.57 24.96 ;
    RECT 55.05 24.2 55.265 24.96 ;
    RECT 55.745 24.2 55.965 24.96 ;
    RECT 56.445 24.2 56.665 24.96 ;
    RECT 57.145 24.2 58.06 24.96 ;
    RECT 58.54 24.2 59.46 24.96 ;
    RECT 59.94 24.2 60.16 24.96 ;
    RECT 60.64 24.2 60.855 24.96 ;
    RECT 61.335 24.2 61.555 24.96 ;
    RECT 62.035 24.2 62.25 24.96 ;
    RECT 62.73 24.2 63.65 24.96 ;
    RECT 64.13 24.2 64.345 24.96 ;
    RECT 64.825 24.2 65.045 24.96 ;
    RECT 65.525 24.2 65.745 24.96 ;
    RECT 66.225 24.2 66.445 24.96 ;
    RECT 66.925 24.2 67.14 24.96 ;
    RECT 67.62 24.2 67.84 24.96 ;
    RECT 68.32 24.2 69.235 24.96 ;
    RECT 69.715 24.2 69.935 24.96 ;
    RECT 70.415 24.2 70.635 24.96 ;
    RECT 71.115 24.2 71.335 24.96 ;
    RECT 71.815 24.2 72.035 24.96 ;
    RECT 72.515 24.2 72.735 24.96 ;
    RECT 73.215 24.2 73.435 24.96 ;
    RECT 73.915 24.2 74.835 24.96 ;
    RECT 75.315 24.2 75.535 24.96 ;
    RECT 76.015 24.2 76.225 24.96 ;
    RECT 76.705 24.2 76.92 24.96 ;
    RECT 77.4 24.2 77.62 24.96 ;
    RECT 78.1 24.2 78.32 24.96 ;
    RECT 78.8 24.2 79.02 24.96 ;
    RECT 79.5 24.2 81.115 24.96 ;
    RECT 81.595 24.2 81.815 24.96 ;
    RECT 82.295 24.2 82.515 24.96 ;
    RECT 82.995 24.2 83.055 24.96 ;
    RECT 83.055 24.11 83.335 25.05 ;
    RECT 83.335 24.2 83.505 24.96 ;
    RECT 26.71 23.44 26.88 24.2 ;
    RECT 26.88 23.35 27.16 24.29 ;
    RECT 27.16 23.44 27.32 24.2 ;
    RECT 27.8 23.44 28.02 24.2 ;
    RECT 28.5 23.44 28.72 24.2 ;
    RECT 29.2 23.44 30.815 24.2 ;
    RECT 31.295 23.44 31.515 24.2 ;
    RECT 31.995 23.44 32.21 24.2 ;
    RECT 32.69 23.44 32.91 24.2 ;
    RECT 33.39 23.44 33.61 24.2 ;
    RECT 34.09 23.44 34.31 24.2 ;
    RECT 34.79 23.44 35.005 24.2 ;
    RECT 35.485 23.44 36.405 24.2 ;
    RECT 36.885 23.44 37.105 24.2 ;
    RECT 37.585 23.44 37.8 24.2 ;
    RECT 38.28 23.44 38.5 24.2 ;
    RECT 38.98 23.44 39.2 24.2 ;
    RECT 39.68 23.44 39.895 24.2 ;
    RECT 40.375 23.44 40.595 24.2 ;
    RECT 41.075 23.44 41.995 24.2 ;
    RECT 42.475 23.44 42.69 24.2 ;
    RECT 43.17 23.44 43.39 24.2 ;
    RECT 43.87 23.44 44.09 24.2 ;
    RECT 44.57 23.44 44.79 24.2 ;
    RECT 45.27 23.44 45.485 24.2 ;
    RECT 45.965 23.44 46.185 24.2 ;
    RECT 46.665 23.44 47.58 24.2 ;
    RECT 48.06 23.44 48.28 24.2 ;
    RECT 48.76 23.44 48.98 24.2 ;
    RECT 49.46 23.44 49.68 24.2 ;
    RECT 50.16 23.44 50.375 24.2 ;
    RECT 50.855 23.44 51.775 24.2 ;
    RECT 52.255 23.44 53.17 24.2 ;
    RECT 53.65 23.44 53.87 24.2 ;
    RECT 54.35 23.44 54.57 24.2 ;
    RECT 55.05 23.44 55.265 24.2 ;
    RECT 55.745 23.44 55.965 24.2 ;
    RECT 56.445 23.44 56.665 24.2 ;
    RECT 57.145 23.44 58.06 24.2 ;
    RECT 58.54 23.44 59.46 24.2 ;
    RECT 59.94 23.44 60.16 24.2 ;
    RECT 60.64 23.44 60.855 24.2 ;
    RECT 61.335 23.44 61.555 24.2 ;
    RECT 62.035 23.44 62.25 24.2 ;
    RECT 62.73 23.44 63.65 24.2 ;
    RECT 64.13 23.44 64.345 24.2 ;
    RECT 64.825 23.44 65.045 24.2 ;
    RECT 65.525 23.44 65.745 24.2 ;
    RECT 66.225 23.44 66.445 24.2 ;
    RECT 66.925 23.44 67.14 24.2 ;
    RECT 67.62 23.44 67.84 24.2 ;
    RECT 68.32 23.44 69.235 24.2 ;
    RECT 69.715 23.44 69.935 24.2 ;
    RECT 70.415 23.44 70.635 24.2 ;
    RECT 71.115 23.44 71.335 24.2 ;
    RECT 71.815 23.44 72.035 24.2 ;
    RECT 72.515 23.44 72.735 24.2 ;
    RECT 73.215 23.44 73.435 24.2 ;
    RECT 73.915 23.44 74.835 24.2 ;
    RECT 75.315 23.44 75.535 24.2 ;
    RECT 76.015 23.44 76.225 24.2 ;
    RECT 76.705 23.44 76.92 24.2 ;
    RECT 77.4 23.44 77.62 24.2 ;
    RECT 78.1 23.44 78.32 24.2 ;
    RECT 78.8 23.44 79.02 24.2 ;
    RECT 79.5 23.44 81.115 24.2 ;
    RECT 81.595 23.44 81.815 24.2 ;
    RECT 82.295 23.44 82.515 24.2 ;
    RECT 82.995 23.44 83.055 24.2 ;
    RECT 83.055 23.35 83.335 24.29 ;
    RECT 83.335 23.44 83.505 24.2 ;
    RECT 4.1 110.77 4.38 110.975 ;
    RECT 7.2 110.77 7.48 110.975 ;
    RECT 10.3 110.77 10.58 110.975 ;
    RECT 13.4 110.77 13.68 110.975 ;
    RECT 16.5 110.77 16.78 110.975 ;
    RECT 19.6 110.77 19.88 110.975 ;
    RECT 22.7 110.77 22.98 110.975 ;
    RECT 1.0 110.77 1.28 110.975 ;
    RECT 19.6 31.8 19.88 32.56 ;
    RECT 19.6 31.04 19.88 31.8 ;
    RECT 19.6 30.28 19.88 31.04 ;
    RECT 19.6 29.52 19.88 30.28 ;
    RECT 19.6 28.76 19.88 29.52 ;
    RECT 19.6 28.0 19.88 28.76 ;
    RECT 19.6 27.24 19.88 28.0 ;
    RECT 19.6 26.48 19.88 27.24 ;
    RECT 19.6 100.18 19.88 100.94 ;
    RECT 19.6 25.72 19.88 26.48 ;
    RECT 19.6 99.42 19.88 100.18 ;
    RECT 19.6 24.96 19.88 25.72 ;
    RECT 19.6 98.66 19.88 99.42 ;
    RECT 19.6 97.9 19.88 98.66 ;
    RECT 19.6 97.14 19.88 97.9 ;
    RECT 19.6 96.38 19.88 97.14 ;
    RECT 19.6 95.62 19.88 96.38 ;
    RECT 19.6 94.86 19.88 95.62 ;
    RECT 19.6 94.1 19.88 94.86 ;
    RECT 19.6 93.34 19.88 94.1 ;
    RECT 19.6 24.2 19.88 24.96 ;
    RECT 19.6 23.44 19.88 24.2 ;
    RECT 19.6 22.68 19.88 23.44 ;
    RECT 19.6 21.92 19.88 22.68 ;
    RECT 19.6 21.16 19.88 21.92 ;
    RECT 19.6 20.4 19.88 21.16 ;
    RECT 19.6 19.64 19.88 20.4 ;
    RECT 19.6 18.88 19.88 19.64 ;
    RECT 19.6 92.58 19.88 93.34 ;
    RECT 19.6 18.12 19.88 18.88 ;
    RECT 19.6 91.82 19.88 92.58 ;
    RECT 19.6 17.36 19.88 18.12 ;
    RECT 19.6 91.06 19.88 91.82 ;
    RECT 19.6 90.3 19.88 91.06 ;
    RECT 19.6 89.54 19.88 90.3 ;
    RECT 19.6 88.78 19.88 89.54 ;
    RECT 19.6 88.02 19.88 88.78 ;
    RECT 19.6 87.26 19.88 88.02 ;
    RECT 19.6 86.5 19.88 87.26 ;
    RECT 19.6 85.74 19.88 86.5 ;
    RECT 19.6 84.98 19.88 85.74 ;
    RECT 19.6 84.22 19.88 84.98 ;
    RECT 19.6 83.46 19.88 84.22 ;
    RECT 19.6 82.7 19.88 83.46 ;
    RECT 19.6 81.94 19.88 82.7 ;
    RECT 19.6 81.18 19.88 81.94 ;
    RECT 19.6 80.42 19.88 81.18 ;
    RECT 19.6 79.66 19.88 80.42 ;
    RECT 19.6 78.9 19.88 79.66 ;
    RECT 19.6 78.14 19.88 78.9 ;
    RECT 19.6 77.38 19.88 78.14 ;
    RECT 19.6 76.62 19.88 77.38 ;
    RECT 19.6 75.86 19.88 76.62 ;
    RECT 19.6 75.1 19.88 75.86 ;
    RECT 19.6 74.34 19.88 75.1 ;
    RECT 19.6 73.58 19.88 74.34 ;
    RECT 19.6 72.82 19.88 73.58 ;
    RECT 19.6 72.06 19.88 72.82 ;
    RECT 19.6 71.3 19.88 72.06 ;
    RECT 19.6 70.54 19.88 71.3 ;
    RECT 19.6 69.78 19.88 70.54 ;
    RECT 19.6 69.02 19.88 69.78 ;
    RECT 19.6 68.26 19.88 69.02 ;
    RECT 19.6 67.5 19.88 68.26 ;
    RECT 19.6 66.74 19.88 67.5 ;
    RECT 19.6 65.98 19.88 66.74 ;
    RECT 19.6 65.22 19.88 65.98 ;
    RECT 19.6 64.46 19.88 65.22 ;
    RECT 19.6 63.7 19.88 64.46 ;
    RECT 19.6 62.94 19.88 63.7 ;
    RECT 19.6 108.54 19.88 109.3 ;
    RECT 19.6 62.18 19.88 62.94 ;
    RECT 19.6 61.42 19.88 62.18 ;
    RECT 19.6 60.66 19.88 61.42 ;
    RECT 19.6 59.92 19.88 60.66 ;
    RECT 19.6 59.16 19.88 59.92 ;
    RECT 19.6 58.4 19.88 59.16 ;
    RECT 19.6 57.64 19.88 58.4 ;
    RECT 19.6 56.88 19.88 57.64 ;
    RECT 19.6 56.12 19.88 56.88 ;
    RECT 19.6 55.36 19.88 56.12 ;
    RECT 19.6 16.6 19.88 17.36 ;
    RECT 19.6 15.84 19.88 16.6 ;
    RECT 19.6 15.08 19.88 15.84 ;
    RECT 19.6 14.32 19.88 15.08 ;
    RECT 19.6 13.56 19.88 14.32 ;
    RECT 19.6 12.8 19.88 13.56 ;
    RECT 19.6 12.04 19.88 12.8 ;
    RECT 19.6 9.81 19.88 11.28 ;
    RECT 19.6 54.6 19.88 55.36 ;
    RECT 19.6 53.84 19.88 54.6 ;
    RECT 19.6 53.08 19.88 53.84 ;
    RECT 19.6 52.32 19.88 53.08 ;
    RECT 19.6 51.56 19.88 52.32 ;
    RECT 19.6 50.8 19.88 51.56 ;
    RECT 19.6 50.04 19.88 50.8 ;
    RECT 19.6 49.28 19.88 50.04 ;
    RECT 19.6 48.52 19.88 49.28 ;
    RECT 19.6 47.76 19.88 48.52 ;
    RECT 19.6 11.28 19.88 12.04 ;
    RECT 19.6 47.0 19.88 47.76 ;
    RECT 19.6 46.24 19.88 47.0 ;
    RECT 19.6 45.48 19.88 46.24 ;
    RECT 19.6 44.72 19.88 45.48 ;
    RECT 19.6 43.96 19.88 44.72 ;
    RECT 19.6 43.2 19.88 43.96 ;
    RECT 19.6 42.44 19.88 43.2 ;
    RECT 19.6 41.68 19.88 42.44 ;
    RECT 19.6 40.92 19.88 41.68 ;
    RECT 19.6 40.16 19.88 40.92 ;
    RECT 19.6 109.3 19.88 110.77 ;
    RECT 19.6 39.4 19.88 40.16 ;
    RECT 19.6 38.64 19.88 39.4 ;
    RECT 19.6 37.88 19.88 38.64 ;
    RECT 19.6 37.12 19.88 37.88 ;
    RECT 19.6 36.36 19.88 37.12 ;
    RECT 19.6 35.6 19.88 36.36 ;
    RECT 19.6 34.84 19.88 35.6 ;
    RECT 19.6 34.08 19.88 34.84 ;
    RECT 19.6 107.78 19.88 108.54 ;
    RECT 19.6 33.32 19.88 34.08 ;
    RECT 19.6 107.02 19.88 107.78 ;
    RECT 19.6 32.56 19.88 33.32 ;
    RECT 19.6 106.26 19.88 107.02 ;
    RECT 19.6 105.5 19.88 106.26 ;
    RECT 19.6 104.74 19.88 105.5 ;
    RECT 19.6 103.98 19.88 104.74 ;
    RECT 19.6 103.22 19.88 103.98 ;
    RECT 19.6 102.46 19.88 103.22 ;
    RECT 19.6 101.7 19.88 102.46 ;
    RECT 19.6 100.94 19.88 101.7 ;
    RECT 7.2 31.8 7.48 32.56 ;
    RECT 7.2 31.04 7.48 31.8 ;
    RECT 7.2 30.28 7.48 31.04 ;
    RECT 7.2 29.52 7.48 30.28 ;
    RECT 7.2 28.76 7.48 29.52 ;
    RECT 7.2 28.0 7.48 28.76 ;
    RECT 7.2 27.24 7.48 28.0 ;
    RECT 7.2 26.48 7.48 27.24 ;
    RECT 7.2 100.18 7.48 100.94 ;
    RECT 7.2 25.72 7.48 26.48 ;
    RECT 7.2 99.42 7.48 100.18 ;
    RECT 7.2 24.96 7.48 25.72 ;
    RECT 7.2 98.66 7.48 99.42 ;
    RECT 7.2 97.9 7.48 98.66 ;
    RECT 7.2 97.14 7.48 97.9 ;
    RECT 7.2 96.38 7.48 97.14 ;
    RECT 7.2 95.62 7.48 96.38 ;
    RECT 7.2 94.86 7.48 95.62 ;
    RECT 7.2 94.1 7.48 94.86 ;
    RECT 7.2 93.34 7.48 94.1 ;
    RECT 7.2 24.2 7.48 24.96 ;
    RECT 7.2 23.44 7.48 24.2 ;
    RECT 7.2 22.68 7.48 23.44 ;
    RECT 7.2 21.92 7.48 22.68 ;
    RECT 7.2 21.16 7.48 21.92 ;
    RECT 7.2 20.4 7.48 21.16 ;
    RECT 7.2 19.64 7.48 20.4 ;
    RECT 7.2 18.88 7.48 19.64 ;
    RECT 7.2 92.58 7.48 93.34 ;
    RECT 7.2 18.12 7.48 18.88 ;
    RECT 7.2 91.82 7.48 92.58 ;
    RECT 7.2 17.36 7.48 18.12 ;
    RECT 7.2 91.06 7.48 91.82 ;
    RECT 7.2 90.3 7.48 91.06 ;
    RECT 7.2 89.54 7.48 90.3 ;
    RECT 7.2 88.78 7.48 89.54 ;
    RECT 7.2 88.02 7.48 88.78 ;
    RECT 7.2 87.26 7.48 88.02 ;
    RECT 7.2 86.5 7.48 87.26 ;
    RECT 7.2 85.74 7.48 86.5 ;
    RECT 7.2 84.98 7.48 85.74 ;
    RECT 7.2 84.22 7.48 84.98 ;
    RECT 7.2 83.46 7.48 84.22 ;
    RECT 7.2 82.7 7.48 83.46 ;
    RECT 7.2 81.94 7.48 82.7 ;
    RECT 7.2 81.18 7.48 81.94 ;
    RECT 7.2 80.42 7.48 81.18 ;
    RECT 7.2 79.66 7.48 80.42 ;
    RECT 7.2 78.9 7.48 79.66 ;
    RECT 7.2 78.14 7.48 78.9 ;
    RECT 7.2 77.38 7.48 78.14 ;
    RECT 7.2 76.62 7.48 77.38 ;
    RECT 7.2 75.86 7.48 76.62 ;
    RECT 7.2 75.1 7.48 75.86 ;
    RECT 7.2 74.34 7.48 75.1 ;
    RECT 7.2 73.58 7.48 74.34 ;
    RECT 7.2 72.82 7.48 73.58 ;
    RECT 7.2 72.06 7.48 72.82 ;
    RECT 7.2 71.3 7.48 72.06 ;
    RECT 7.2 70.54 7.48 71.3 ;
    RECT 7.2 69.78 7.48 70.54 ;
    RECT 7.2 69.02 7.48 69.78 ;
    RECT 7.2 68.26 7.48 69.02 ;
    RECT 7.2 67.5 7.48 68.26 ;
    RECT 7.2 66.74 7.48 67.5 ;
    RECT 7.2 65.98 7.48 66.74 ;
    RECT 7.2 65.22 7.48 65.98 ;
    RECT 7.2 64.46 7.48 65.22 ;
    RECT 7.2 63.7 7.48 64.46 ;
    RECT 7.2 62.94 7.48 63.7 ;
    RECT 7.2 108.54 7.48 109.3 ;
    RECT 7.2 62.18 7.48 62.94 ;
    RECT 7.2 61.42 7.48 62.18 ;
    RECT 7.2 60.66 7.48 61.42 ;
    RECT 7.2 59.92 7.48 60.66 ;
    RECT 7.2 59.16 7.48 59.92 ;
    RECT 7.2 58.4 7.48 59.16 ;
    RECT 7.2 57.64 7.48 58.4 ;
    RECT 7.2 56.88 7.48 57.64 ;
    RECT 7.2 56.12 7.48 56.88 ;
    RECT 7.2 55.36 7.48 56.12 ;
    RECT 7.2 16.6 7.48 17.36 ;
    RECT 7.2 15.84 7.48 16.6 ;
    RECT 7.2 15.08 7.48 15.84 ;
    RECT 7.2 14.32 7.48 15.08 ;
    RECT 7.2 13.56 7.48 14.32 ;
    RECT 7.2 12.8 7.48 13.56 ;
    RECT 7.2 12.04 7.48 12.8 ;
    RECT 7.2 9.81 7.48 11.28 ;
    RECT 7.2 54.6 7.48 55.36 ;
    RECT 7.2 53.84 7.48 54.6 ;
    RECT 7.2 53.08 7.48 53.84 ;
    RECT 7.2 52.32 7.48 53.08 ;
    RECT 7.2 51.56 7.48 52.32 ;
    RECT 7.2 50.8 7.48 51.56 ;
    RECT 7.2 50.04 7.48 50.8 ;
    RECT 7.2 49.28 7.48 50.04 ;
    RECT 7.2 48.52 7.48 49.28 ;
    RECT 7.2 47.76 7.48 48.52 ;
    RECT 7.2 11.28 7.48 12.04 ;
    RECT 7.2 47.0 7.48 47.76 ;
    RECT 7.2 46.24 7.48 47.0 ;
    RECT 7.2 45.48 7.48 46.24 ;
    RECT 7.2 44.72 7.48 45.48 ;
    RECT 7.2 43.96 7.48 44.72 ;
    RECT 7.2 43.2 7.48 43.96 ;
    RECT 7.2 42.44 7.48 43.2 ;
    RECT 7.2 41.68 7.48 42.44 ;
    RECT 7.2 40.92 7.48 41.68 ;
    RECT 7.2 40.16 7.48 40.92 ;
    RECT 7.2 109.3 7.48 110.77 ;
    RECT 7.2 39.4 7.48 40.16 ;
    RECT 7.2 38.64 7.48 39.4 ;
    RECT 7.2 37.88 7.48 38.64 ;
    RECT 7.2 37.12 7.48 37.88 ;
    RECT 7.2 36.36 7.48 37.12 ;
    RECT 7.2 35.6 7.48 36.36 ;
    RECT 7.2 34.84 7.48 35.6 ;
    RECT 7.2 34.08 7.48 34.84 ;
    RECT 7.2 107.78 7.48 108.54 ;
    RECT 7.2 33.32 7.48 34.08 ;
    RECT 7.2 107.02 7.48 107.78 ;
    RECT 7.2 32.56 7.48 33.32 ;
    RECT 7.2 106.26 7.48 107.02 ;
    RECT 7.2 105.5 7.48 106.26 ;
    RECT 7.2 104.74 7.48 105.5 ;
    RECT 7.2 103.98 7.48 104.74 ;
    RECT 7.2 103.22 7.48 103.98 ;
    RECT 7.2 102.46 7.48 103.22 ;
    RECT 7.2 101.7 7.48 102.46 ;
    RECT 7.2 100.94 7.48 101.7 ;
    RECT 10.3 31.8 10.58 32.56 ;
    RECT 10.3 31.04 10.58 31.8 ;
    RECT 10.3 30.28 10.58 31.04 ;
    RECT 10.3 29.52 10.58 30.28 ;
    RECT 10.3 28.76 10.58 29.52 ;
    RECT 10.3 28.0 10.58 28.76 ;
    RECT 10.3 27.24 10.58 28.0 ;
    RECT 10.3 26.48 10.58 27.24 ;
    RECT 10.3 100.18 10.58 100.94 ;
    RECT 10.3 25.72 10.58 26.48 ;
    RECT 10.3 99.42 10.58 100.18 ;
    RECT 10.3 24.96 10.58 25.72 ;
    RECT 10.3 98.66 10.58 99.42 ;
    RECT 10.3 97.9 10.58 98.66 ;
    RECT 10.3 97.14 10.58 97.9 ;
    RECT 10.3 96.38 10.58 97.14 ;
    RECT 10.3 95.62 10.58 96.38 ;
    RECT 10.3 94.86 10.58 95.62 ;
    RECT 10.3 94.1 10.58 94.86 ;
    RECT 10.3 93.34 10.58 94.1 ;
    RECT 10.3 24.2 10.58 24.96 ;
    RECT 10.3 23.44 10.58 24.2 ;
    RECT 10.3 22.68 10.58 23.44 ;
    RECT 10.3 21.92 10.58 22.68 ;
    RECT 10.3 21.16 10.58 21.92 ;
    RECT 10.3 20.4 10.58 21.16 ;
    RECT 10.3 19.64 10.58 20.4 ;
    RECT 10.3 18.88 10.58 19.64 ;
    RECT 10.3 92.58 10.58 93.34 ;
    RECT 10.3 18.12 10.58 18.88 ;
    RECT 10.3 91.82 10.58 92.58 ;
    RECT 10.3 17.36 10.58 18.12 ;
    RECT 10.3 91.06 10.58 91.82 ;
    RECT 10.3 90.3 10.58 91.06 ;
    RECT 10.3 89.54 10.58 90.3 ;
    RECT 10.3 88.78 10.58 89.54 ;
    RECT 10.3 88.02 10.58 88.78 ;
    RECT 10.3 87.26 10.58 88.02 ;
    RECT 10.3 86.5 10.58 87.26 ;
    RECT 10.3 85.74 10.58 86.5 ;
    RECT 10.3 84.98 10.58 85.74 ;
    RECT 10.3 84.22 10.58 84.98 ;
    RECT 10.3 83.46 10.58 84.22 ;
    RECT 10.3 82.7 10.58 83.46 ;
    RECT 10.3 81.94 10.58 82.7 ;
    RECT 10.3 81.18 10.58 81.94 ;
    RECT 10.3 80.42 10.58 81.18 ;
    RECT 10.3 79.66 10.58 80.42 ;
    RECT 10.3 78.9 10.58 79.66 ;
    RECT 10.3 78.14 10.58 78.9 ;
    RECT 10.3 77.38 10.58 78.14 ;
    RECT 10.3 76.62 10.58 77.38 ;
    RECT 10.3 75.86 10.58 76.62 ;
    RECT 10.3 75.1 10.58 75.86 ;
    RECT 10.3 74.34 10.58 75.1 ;
    RECT 10.3 73.58 10.58 74.34 ;
    RECT 10.3 72.82 10.58 73.58 ;
    RECT 10.3 72.06 10.58 72.82 ;
    RECT 10.3 71.3 10.58 72.06 ;
    RECT 10.3 70.54 10.58 71.3 ;
    RECT 10.3 69.78 10.58 70.54 ;
    RECT 10.3 69.02 10.58 69.78 ;
    RECT 10.3 68.26 10.58 69.02 ;
    RECT 10.3 67.5 10.58 68.26 ;
    RECT 10.3 66.74 10.58 67.5 ;
    RECT 10.3 65.98 10.58 66.74 ;
    RECT 10.3 65.22 10.58 65.98 ;
    RECT 10.3 64.46 10.58 65.22 ;
    RECT 10.3 63.7 10.58 64.46 ;
    RECT 10.3 62.94 10.58 63.7 ;
    RECT 10.3 108.54 10.58 109.3 ;
    RECT 10.3 62.18 10.58 62.94 ;
    RECT 10.3 61.42 10.58 62.18 ;
    RECT 10.3 60.66 10.58 61.42 ;
    RECT 10.3 59.92 10.58 60.66 ;
    RECT 10.3 59.16 10.58 59.92 ;
    RECT 10.3 58.4 10.58 59.16 ;
    RECT 10.3 57.64 10.58 58.4 ;
    RECT 10.3 56.88 10.58 57.64 ;
    RECT 10.3 56.12 10.58 56.88 ;
    RECT 10.3 55.36 10.58 56.12 ;
    RECT 10.3 16.6 10.58 17.36 ;
    RECT 10.3 15.84 10.58 16.6 ;
    RECT 10.3 15.08 10.58 15.84 ;
    RECT 10.3 14.32 10.58 15.08 ;
    RECT 10.3 13.56 10.58 14.32 ;
    RECT 10.3 12.8 10.58 13.56 ;
    RECT 10.3 12.04 10.58 12.8 ;
    RECT 10.3 9.81 10.58 11.28 ;
    RECT 10.3 54.6 10.58 55.36 ;
    RECT 10.3 53.84 10.58 54.6 ;
    RECT 10.3 53.08 10.58 53.84 ;
    RECT 10.3 52.32 10.58 53.08 ;
    RECT 10.3 51.56 10.58 52.32 ;
    RECT 10.3 50.8 10.58 51.56 ;
    RECT 10.3 50.04 10.58 50.8 ;
    RECT 10.3 49.28 10.58 50.04 ;
    RECT 10.3 48.52 10.58 49.28 ;
    RECT 10.3 47.76 10.58 48.52 ;
    RECT 10.3 11.28 10.58 12.04 ;
    RECT 10.3 47.0 10.58 47.76 ;
    RECT 10.3 46.24 10.58 47.0 ;
    RECT 10.3 45.48 10.58 46.24 ;
    RECT 10.3 44.72 10.58 45.48 ;
    RECT 10.3 43.96 10.58 44.72 ;
    RECT 10.3 43.2 10.58 43.96 ;
    RECT 10.3 42.44 10.58 43.2 ;
    RECT 10.3 41.68 10.58 42.44 ;
    RECT 10.3 40.92 10.58 41.68 ;
    RECT 10.3 40.16 10.58 40.92 ;
    RECT 10.3 109.3 10.58 110.77 ;
    RECT 10.3 39.4 10.58 40.16 ;
    RECT 10.3 38.64 10.58 39.4 ;
    RECT 10.3 37.88 10.58 38.64 ;
    RECT 10.3 37.12 10.58 37.88 ;
    RECT 10.3 36.36 10.58 37.12 ;
    RECT 10.3 35.6 10.58 36.36 ;
    RECT 10.3 34.84 10.58 35.6 ;
    RECT 10.3 34.08 10.58 34.84 ;
    RECT 10.3 107.78 10.58 108.54 ;
    RECT 10.3 33.32 10.58 34.08 ;
    RECT 10.3 107.02 10.58 107.78 ;
    RECT 10.3 32.56 10.58 33.32 ;
    RECT 10.3 106.26 10.58 107.02 ;
    RECT 10.3 105.5 10.58 106.26 ;
    RECT 10.3 104.74 10.58 105.5 ;
    RECT 10.3 103.98 10.58 104.74 ;
    RECT 10.3 103.22 10.58 103.98 ;
    RECT 10.3 102.46 10.58 103.22 ;
    RECT 10.3 101.7 10.58 102.46 ;
    RECT 10.3 100.94 10.58 101.7 ;
    RECT 13.4 31.8 13.68 32.56 ;
    RECT 13.4 31.04 13.68 31.8 ;
    RECT 13.4 30.28 13.68 31.04 ;
    RECT 13.4 29.52 13.68 30.28 ;
    RECT 13.4 28.76 13.68 29.52 ;
    RECT 13.4 28.0 13.68 28.76 ;
    RECT 13.4 27.24 13.68 28.0 ;
    RECT 13.4 26.48 13.68 27.24 ;
    RECT 13.4 100.18 13.68 100.94 ;
    RECT 13.4 25.72 13.68 26.48 ;
    RECT 13.4 99.42 13.68 100.18 ;
    RECT 13.4 24.96 13.68 25.72 ;
    RECT 13.4 98.66 13.68 99.42 ;
    RECT 13.4 97.9 13.68 98.66 ;
    RECT 13.4 97.14 13.68 97.9 ;
    RECT 13.4 96.38 13.68 97.14 ;
    RECT 13.4 95.62 13.68 96.38 ;
    RECT 13.4 94.86 13.68 95.62 ;
    RECT 13.4 94.1 13.68 94.86 ;
    RECT 13.4 93.34 13.68 94.1 ;
    RECT 13.4 24.2 13.68 24.96 ;
    RECT 13.4 23.44 13.68 24.2 ;
    RECT 13.4 22.68 13.68 23.44 ;
    RECT 13.4 21.92 13.68 22.68 ;
    RECT 13.4 21.16 13.68 21.92 ;
    RECT 13.4 20.4 13.68 21.16 ;
    RECT 13.4 19.64 13.68 20.4 ;
    RECT 13.4 18.88 13.68 19.64 ;
    RECT 13.4 92.58 13.68 93.34 ;
    RECT 13.4 18.12 13.68 18.88 ;
    RECT 13.4 91.82 13.68 92.58 ;
    RECT 13.4 17.36 13.68 18.12 ;
    RECT 13.4 91.06 13.68 91.82 ;
    RECT 13.4 90.3 13.68 91.06 ;
    RECT 13.4 89.54 13.68 90.3 ;
    RECT 13.4 88.78 13.68 89.54 ;
    RECT 13.4 88.02 13.68 88.78 ;
    RECT 13.4 87.26 13.68 88.02 ;
    RECT 13.4 86.5 13.68 87.26 ;
    RECT 13.4 85.74 13.68 86.5 ;
    RECT 13.4 84.98 13.68 85.74 ;
    RECT 13.4 84.22 13.68 84.98 ;
    RECT 13.4 83.46 13.68 84.22 ;
    RECT 13.4 82.7 13.68 83.46 ;
    RECT 13.4 81.94 13.68 82.7 ;
    RECT 13.4 81.18 13.68 81.94 ;
    RECT 13.4 80.42 13.68 81.18 ;
    RECT 13.4 79.66 13.68 80.42 ;
    RECT 13.4 78.9 13.68 79.66 ;
    RECT 13.4 78.14 13.68 78.9 ;
    RECT 13.4 77.38 13.68 78.14 ;
    RECT 13.4 76.62 13.68 77.38 ;
    RECT 13.4 75.86 13.68 76.62 ;
    RECT 13.4 75.1 13.68 75.86 ;
    RECT 13.4 74.34 13.68 75.1 ;
    RECT 13.4 73.58 13.68 74.34 ;
    RECT 13.4 72.82 13.68 73.58 ;
    RECT 13.4 72.06 13.68 72.82 ;
    RECT 13.4 71.3 13.68 72.06 ;
    RECT 13.4 70.54 13.68 71.3 ;
    RECT 13.4 69.78 13.68 70.54 ;
    RECT 13.4 69.02 13.68 69.78 ;
    RECT 13.4 68.26 13.68 69.02 ;
    RECT 13.4 67.5 13.68 68.26 ;
    RECT 13.4 66.74 13.68 67.5 ;
    RECT 13.4 65.98 13.68 66.74 ;
    RECT 13.4 65.22 13.68 65.98 ;
    RECT 13.4 64.46 13.68 65.22 ;
    RECT 13.4 63.7 13.68 64.46 ;
    RECT 13.4 62.94 13.68 63.7 ;
    RECT 13.4 108.54 13.68 109.3 ;
    RECT 13.4 62.18 13.68 62.94 ;
    RECT 13.4 61.42 13.68 62.18 ;
    RECT 13.4 60.66 13.68 61.42 ;
    RECT 13.4 59.92 13.68 60.66 ;
    RECT 13.4 59.16 13.68 59.92 ;
    RECT 13.4 58.4 13.68 59.16 ;
    RECT 13.4 57.64 13.68 58.4 ;
    RECT 13.4 56.88 13.68 57.64 ;
    RECT 13.4 56.12 13.68 56.88 ;
    RECT 13.4 55.36 13.68 56.12 ;
    RECT 13.4 16.6 13.68 17.36 ;
    RECT 13.4 15.84 13.68 16.6 ;
    RECT 13.4 15.08 13.68 15.84 ;
    RECT 13.4 14.32 13.68 15.08 ;
    RECT 13.4 13.56 13.68 14.32 ;
    RECT 13.4 12.8 13.68 13.56 ;
    RECT 13.4 12.04 13.68 12.8 ;
    RECT 13.4 9.81 13.68 11.28 ;
    RECT 13.4 54.6 13.68 55.36 ;
    RECT 13.4 53.84 13.68 54.6 ;
    RECT 13.4 53.08 13.68 53.84 ;
    RECT 13.4 52.32 13.68 53.08 ;
    RECT 13.4 51.56 13.68 52.32 ;
    RECT 13.4 50.8 13.68 51.56 ;
    RECT 13.4 50.04 13.68 50.8 ;
    RECT 13.4 49.28 13.68 50.04 ;
    RECT 13.4 48.52 13.68 49.28 ;
    RECT 13.4 47.76 13.68 48.52 ;
    RECT 13.4 11.28 13.68 12.04 ;
    RECT 13.4 47.0 13.68 47.76 ;
    RECT 13.4 46.24 13.68 47.0 ;
    RECT 13.4 45.48 13.68 46.24 ;
    RECT 13.4 44.72 13.68 45.48 ;
    RECT 13.4 43.96 13.68 44.72 ;
    RECT 13.4 43.2 13.68 43.96 ;
    RECT 13.4 42.44 13.68 43.2 ;
    RECT 13.4 41.68 13.68 42.44 ;
    RECT 13.4 40.92 13.68 41.68 ;
    RECT 13.4 40.16 13.68 40.92 ;
    RECT 13.4 109.3 13.68 110.77 ;
    RECT 13.4 39.4 13.68 40.16 ;
    RECT 13.4 38.64 13.68 39.4 ;
    RECT 13.4 37.88 13.68 38.64 ;
    RECT 13.4 37.12 13.68 37.88 ;
    RECT 13.4 36.36 13.68 37.12 ;
    RECT 13.4 35.6 13.68 36.36 ;
    RECT 13.4 34.84 13.68 35.6 ;
    RECT 13.4 34.08 13.68 34.84 ;
    RECT 13.4 107.78 13.68 108.54 ;
    RECT 13.4 33.32 13.68 34.08 ;
    RECT 13.4 107.02 13.68 107.78 ;
    RECT 13.4 32.56 13.68 33.32 ;
    RECT 13.4 106.26 13.68 107.02 ;
    RECT 13.4 105.5 13.68 106.26 ;
    RECT 13.4 104.74 13.68 105.5 ;
    RECT 13.4 103.98 13.68 104.74 ;
    RECT 13.4 103.22 13.68 103.98 ;
    RECT 13.4 102.46 13.68 103.22 ;
    RECT 13.4 101.7 13.68 102.46 ;
    RECT 13.4 100.94 13.68 101.7 ;
    RECT 16.5 31.8 16.78 32.56 ;
    RECT 16.5 31.04 16.78 31.8 ;
    RECT 16.5 30.28 16.78 31.04 ;
    RECT 16.5 29.52 16.78 30.28 ;
    RECT 16.5 28.76 16.78 29.52 ;
    RECT 16.5 28.0 16.78 28.76 ;
    RECT 16.5 27.24 16.78 28.0 ;
    RECT 16.5 26.48 16.78 27.24 ;
    RECT 16.5 100.18 16.78 100.94 ;
    RECT 16.5 25.72 16.78 26.48 ;
    RECT 16.5 99.42 16.78 100.18 ;
    RECT 16.5 24.96 16.78 25.72 ;
    RECT 16.5 98.66 16.78 99.42 ;
    RECT 16.5 97.9 16.78 98.66 ;
    RECT 16.5 97.14 16.78 97.9 ;
    RECT 16.5 96.38 16.78 97.14 ;
    RECT 16.5 95.62 16.78 96.38 ;
    RECT 16.5 94.86 16.78 95.62 ;
    RECT 16.5 94.1 16.78 94.86 ;
    RECT 16.5 93.34 16.78 94.1 ;
    RECT 16.5 24.2 16.78 24.96 ;
    RECT 16.5 23.44 16.78 24.2 ;
    RECT 16.5 22.68 16.78 23.44 ;
    RECT 16.5 21.92 16.78 22.68 ;
    RECT 16.5 21.16 16.78 21.92 ;
    RECT 16.5 20.4 16.78 21.16 ;
    RECT 16.5 19.64 16.78 20.4 ;
    RECT 16.5 18.88 16.78 19.64 ;
    RECT 16.5 92.58 16.78 93.34 ;
    RECT 16.5 18.12 16.78 18.88 ;
    RECT 16.5 91.82 16.78 92.58 ;
    RECT 16.5 17.36 16.78 18.12 ;
    RECT 16.5 91.06 16.78 91.82 ;
    RECT 16.5 90.3 16.78 91.06 ;
    RECT 16.5 89.54 16.78 90.3 ;
    RECT 16.5 88.78 16.78 89.54 ;
    RECT 16.5 88.02 16.78 88.78 ;
    RECT 16.5 87.26 16.78 88.02 ;
    RECT 16.5 86.5 16.78 87.26 ;
    RECT 16.5 85.74 16.78 86.5 ;
    RECT 16.5 84.98 16.78 85.74 ;
    RECT 16.5 84.22 16.78 84.98 ;
    RECT 16.5 83.46 16.78 84.22 ;
    RECT 16.5 82.7 16.78 83.46 ;
    RECT 16.5 81.94 16.78 82.7 ;
    RECT 16.5 81.18 16.78 81.94 ;
    RECT 16.5 80.42 16.78 81.18 ;
    RECT 16.5 79.66 16.78 80.42 ;
    RECT 16.5 78.9 16.78 79.66 ;
    RECT 16.5 78.14 16.78 78.9 ;
    RECT 16.5 77.38 16.78 78.14 ;
    RECT 16.5 76.62 16.78 77.38 ;
    RECT 16.5 75.86 16.78 76.62 ;
    RECT 16.5 75.1 16.78 75.86 ;
    RECT 16.5 74.34 16.78 75.1 ;
    RECT 16.5 73.58 16.78 74.34 ;
    RECT 16.5 72.82 16.78 73.58 ;
    RECT 16.5 72.06 16.78 72.82 ;
    RECT 16.5 71.3 16.78 72.06 ;
    RECT 16.5 70.54 16.78 71.3 ;
    RECT 16.5 69.78 16.78 70.54 ;
    RECT 16.5 69.02 16.78 69.78 ;
    RECT 16.5 68.26 16.78 69.02 ;
    RECT 16.5 67.5 16.78 68.26 ;
    RECT 16.5 66.74 16.78 67.5 ;
    RECT 16.5 65.98 16.78 66.74 ;
    RECT 16.5 65.22 16.78 65.98 ;
    RECT 16.5 64.46 16.78 65.22 ;
    RECT 16.5 63.7 16.78 64.46 ;
    RECT 16.5 62.94 16.78 63.7 ;
    RECT 16.5 108.54 16.78 109.3 ;
    RECT 16.5 62.18 16.78 62.94 ;
    RECT 16.5 61.42 16.78 62.18 ;
    RECT 16.5 60.66 16.78 61.42 ;
    RECT 16.5 59.92 16.78 60.66 ;
    RECT 16.5 59.16 16.78 59.92 ;
    RECT 16.5 58.4 16.78 59.16 ;
    RECT 16.5 57.64 16.78 58.4 ;
    RECT 16.5 56.88 16.78 57.64 ;
    RECT 16.5 56.12 16.78 56.88 ;
    RECT 16.5 55.36 16.78 56.12 ;
    RECT 16.5 16.6 16.78 17.36 ;
    RECT 16.5 15.84 16.78 16.6 ;
    RECT 16.5 15.08 16.78 15.84 ;
    RECT 16.5 14.32 16.78 15.08 ;
    RECT 16.5 13.56 16.78 14.32 ;
    RECT 16.5 12.8 16.78 13.56 ;
    RECT 16.5 12.04 16.78 12.8 ;
    RECT 16.5 9.81 16.78 11.28 ;
    RECT 16.5 54.6 16.78 55.36 ;
    RECT 16.5 53.84 16.78 54.6 ;
    RECT 16.5 53.08 16.78 53.84 ;
    RECT 16.5 52.32 16.78 53.08 ;
    RECT 16.5 51.56 16.78 52.32 ;
    RECT 16.5 50.8 16.78 51.56 ;
    RECT 16.5 50.04 16.78 50.8 ;
    RECT 16.5 49.28 16.78 50.04 ;
    RECT 16.5 48.52 16.78 49.28 ;
    RECT 16.5 47.76 16.78 48.52 ;
    RECT 16.5 11.28 16.78 12.04 ;
    RECT 16.5 47.0 16.78 47.76 ;
    RECT 16.5 46.24 16.78 47.0 ;
    RECT 16.5 45.48 16.78 46.24 ;
    RECT 16.5 44.72 16.78 45.48 ;
    RECT 16.5 43.96 16.78 44.72 ;
    RECT 16.5 43.2 16.78 43.96 ;
    RECT 16.5 42.44 16.78 43.2 ;
    RECT 16.5 41.68 16.78 42.44 ;
    RECT 16.5 40.92 16.78 41.68 ;
    RECT 16.5 40.16 16.78 40.92 ;
    RECT 16.5 109.3 16.78 110.77 ;
    RECT 16.5 39.4 16.78 40.16 ;
    RECT 16.5 38.64 16.78 39.4 ;
    RECT 16.5 37.88 16.78 38.64 ;
    RECT 16.5 37.12 16.78 37.88 ;
    RECT 16.5 36.36 16.78 37.12 ;
    RECT 16.5 35.6 16.78 36.36 ;
    RECT 16.5 34.84 16.78 35.6 ;
    RECT 16.5 34.08 16.78 34.84 ;
    RECT 16.5 107.78 16.78 108.54 ;
    RECT 16.5 33.32 16.78 34.08 ;
    RECT 16.5 107.02 16.78 107.78 ;
    RECT 16.5 32.56 16.78 33.32 ;
    RECT 16.5 106.26 16.78 107.02 ;
    RECT 16.5 105.5 16.78 106.26 ;
    RECT 16.5 104.74 16.78 105.5 ;
    RECT 16.5 103.98 16.78 104.74 ;
    RECT 16.5 103.22 16.78 103.98 ;
    RECT 16.5 102.46 16.78 103.22 ;
    RECT 16.5 101.7 16.78 102.46 ;
    RECT 16.5 100.94 16.78 101.7 ;
    RECT 4.1 31.8 4.38 32.56 ;
    RECT 4.1 31.04 4.38 31.8 ;
    RECT 4.1 30.28 4.38 31.04 ;
    RECT 4.1 29.52 4.38 30.28 ;
    RECT 4.1 28.76 4.38 29.52 ;
    RECT 4.1 28.0 4.38 28.76 ;
    RECT 4.1 27.24 4.38 28.0 ;
    RECT 4.1 26.48 4.38 27.24 ;
    RECT 4.1 100.18 4.38 100.94 ;
    RECT 4.1 25.72 4.38 26.48 ;
    RECT 4.1 99.42 4.38 100.18 ;
    RECT 4.1 24.96 4.38 25.72 ;
    RECT 4.1 98.66 4.38 99.42 ;
    RECT 4.1 97.9 4.38 98.66 ;
    RECT 4.1 97.14 4.38 97.9 ;
    RECT 4.1 96.38 4.38 97.14 ;
    RECT 4.1 95.62 4.38 96.38 ;
    RECT 4.1 94.86 4.38 95.62 ;
    RECT 4.1 94.1 4.38 94.86 ;
    RECT 4.1 93.34 4.38 94.1 ;
    RECT 4.1 24.2 4.38 24.96 ;
    RECT 4.1 23.44 4.38 24.2 ;
    RECT 4.1 22.68 4.38 23.44 ;
    RECT 4.1 21.92 4.38 22.68 ;
    RECT 4.1 21.16 4.38 21.92 ;
    RECT 4.1 20.4 4.38 21.16 ;
    RECT 4.1 19.64 4.38 20.4 ;
    RECT 4.1 18.88 4.38 19.64 ;
    RECT 4.1 92.58 4.38 93.34 ;
    RECT 4.1 18.12 4.38 18.88 ;
    RECT 4.1 91.82 4.38 92.58 ;
    RECT 4.1 17.36 4.38 18.12 ;
    RECT 4.1 91.06 4.38 91.82 ;
    RECT 4.1 90.3 4.38 91.06 ;
    RECT 4.1 89.54 4.38 90.3 ;
    RECT 4.1 88.78 4.38 89.54 ;
    RECT 4.1 88.02 4.38 88.78 ;
    RECT 4.1 87.26 4.38 88.02 ;
    RECT 4.1 86.5 4.38 87.26 ;
    RECT 4.1 85.74 4.38 86.5 ;
    RECT 4.1 84.98 4.38 85.74 ;
    RECT 4.1 84.22 4.38 84.98 ;
    RECT 4.1 83.46 4.38 84.22 ;
    RECT 4.1 82.7 4.38 83.46 ;
    RECT 4.1 81.94 4.38 82.7 ;
    RECT 4.1 81.18 4.38 81.94 ;
    RECT 4.1 80.42 4.38 81.18 ;
    RECT 4.1 79.66 4.38 80.42 ;
    RECT 4.1 78.9 4.38 79.66 ;
    RECT 4.1 78.14 4.38 78.9 ;
    RECT 4.1 77.38 4.38 78.14 ;
    RECT 4.1 76.62 4.38 77.38 ;
    RECT 4.1 75.86 4.38 76.62 ;
    RECT 4.1 75.1 4.38 75.86 ;
    RECT 4.1 74.34 4.38 75.1 ;
    RECT 4.1 73.58 4.38 74.34 ;
    RECT 4.1 72.82 4.38 73.58 ;
    RECT 4.1 72.06 4.38 72.82 ;
    RECT 4.1 71.3 4.38 72.06 ;
    RECT 4.1 70.54 4.38 71.3 ;
    RECT 4.1 69.78 4.38 70.54 ;
    RECT 4.1 69.02 4.38 69.78 ;
    RECT 4.1 68.26 4.38 69.02 ;
    RECT 4.1 67.5 4.38 68.26 ;
    RECT 4.1 66.74 4.38 67.5 ;
    RECT 4.1 65.98 4.38 66.74 ;
    RECT 4.1 65.22 4.38 65.98 ;
    RECT 4.1 64.46 4.38 65.22 ;
    RECT 4.1 63.7 4.38 64.46 ;
    RECT 4.1 62.94 4.38 63.7 ;
    RECT 4.1 108.54 4.38 109.3 ;
    RECT 4.1 62.18 4.38 62.94 ;
    RECT 4.1 61.42 4.38 62.18 ;
    RECT 4.1 60.66 4.38 61.42 ;
    RECT 4.1 59.92 4.38 60.66 ;
    RECT 4.1 59.16 4.38 59.92 ;
    RECT 4.1 58.4 4.38 59.16 ;
    RECT 4.1 57.64 4.38 58.4 ;
    RECT 4.1 56.88 4.38 57.64 ;
    RECT 4.1 56.12 4.38 56.88 ;
    RECT 4.1 55.36 4.38 56.12 ;
    RECT 4.1 16.6 4.38 17.36 ;
    RECT 4.1 15.84 4.38 16.6 ;
    RECT 4.1 15.08 4.38 15.84 ;
    RECT 4.1 14.32 4.38 15.08 ;
    RECT 4.1 13.56 4.38 14.32 ;
    RECT 4.1 12.8 4.38 13.56 ;
    RECT 4.1 12.04 4.38 12.8 ;
    RECT 4.1 9.81 4.38 11.28 ;
    RECT 4.1 54.6 4.38 55.36 ;
    RECT 4.1 53.84 4.38 54.6 ;
    RECT 4.1 53.08 4.38 53.84 ;
    RECT 4.1 52.32 4.38 53.08 ;
    RECT 4.1 51.56 4.38 52.32 ;
    RECT 4.1 50.8 4.38 51.56 ;
    RECT 4.1 50.04 4.38 50.8 ;
    RECT 4.1 49.28 4.38 50.04 ;
    RECT 4.1 48.52 4.38 49.28 ;
    RECT 4.1 47.76 4.38 48.52 ;
    RECT 4.1 11.28 4.38 12.04 ;
    RECT 4.1 47.0 4.38 47.76 ;
    RECT 4.1 46.24 4.38 47.0 ;
    RECT 4.1 45.48 4.38 46.24 ;
    RECT 4.1 44.72 4.38 45.48 ;
    RECT 4.1 43.96 4.38 44.72 ;
    RECT 4.1 43.2 4.38 43.96 ;
    RECT 4.1 42.44 4.38 43.2 ;
    RECT 4.1 41.68 4.38 42.44 ;
    RECT 4.1 40.92 4.38 41.68 ;
    RECT 4.1 40.16 4.38 40.92 ;
    RECT 4.1 109.3 4.38 110.77 ;
    RECT 4.1 39.4 4.38 40.16 ;
    RECT 4.1 38.64 4.38 39.4 ;
    RECT 4.1 37.88 4.38 38.64 ;
    RECT 4.1 37.12 4.38 37.88 ;
    RECT 4.1 36.36 4.38 37.12 ;
    RECT 4.1 35.6 4.38 36.36 ;
    RECT 4.1 34.84 4.38 35.6 ;
    RECT 4.1 34.08 4.38 34.84 ;
    RECT 4.1 107.78 4.38 108.54 ;
    RECT 4.1 33.32 4.38 34.08 ;
    RECT 4.1 107.02 4.38 107.78 ;
    RECT 4.1 32.56 4.38 33.32 ;
    RECT 4.1 106.26 4.38 107.02 ;
    RECT 4.1 105.5 4.38 106.26 ;
    RECT 4.1 104.74 4.38 105.5 ;
    RECT 4.1 103.98 4.38 104.74 ;
    RECT 4.1 103.22 4.38 103.98 ;
    RECT 4.1 102.46 4.38 103.22 ;
    RECT 4.1 101.7 4.38 102.46 ;
    RECT 4.1 100.94 4.38 101.7 ;
    RECT 22.7 31.8 22.98 32.56 ;
    RECT 22.7 31.04 22.98 31.8 ;
    RECT 22.7 30.28 22.98 31.04 ;
    RECT 22.7 29.52 22.98 30.28 ;
    RECT 22.7 28.76 22.98 29.52 ;
    RECT 22.7 28.0 22.98 28.76 ;
    RECT 22.7 27.24 22.98 28.0 ;
    RECT 22.7 26.48 22.98 27.24 ;
    RECT 22.7 100.18 22.98 100.94 ;
    RECT 22.7 25.72 22.98 26.48 ;
    RECT 22.7 99.42 22.98 100.18 ;
    RECT 22.7 24.96 22.98 25.72 ;
    RECT 22.7 98.66 22.98 99.42 ;
    RECT 22.7 97.9 22.98 98.66 ;
    RECT 22.7 97.14 22.98 97.9 ;
    RECT 22.7 96.38 22.98 97.14 ;
    RECT 22.7 95.62 22.98 96.38 ;
    RECT 22.7 94.86 22.98 95.62 ;
    RECT 22.7 94.1 22.98 94.86 ;
    RECT 22.7 93.34 22.98 94.1 ;
    RECT 22.7 24.2 22.98 24.96 ;
    RECT 22.7 23.44 22.98 24.2 ;
    RECT 22.7 22.68 22.98 23.44 ;
    RECT 22.7 21.92 22.98 22.68 ;
    RECT 22.7 21.16 22.98 21.92 ;
    RECT 22.7 20.4 22.98 21.16 ;
    RECT 22.7 19.64 22.98 20.4 ;
    RECT 22.7 18.88 22.98 19.64 ;
    RECT 22.7 92.58 22.98 93.34 ;
    RECT 22.7 18.12 22.98 18.88 ;
    RECT 22.7 91.82 22.98 92.58 ;
    RECT 22.7 17.36 22.98 18.12 ;
    RECT 22.7 91.06 22.98 91.82 ;
    RECT 22.7 90.3 22.98 91.06 ;
    RECT 22.7 89.54 22.98 90.3 ;
    RECT 22.7 88.78 22.98 89.54 ;
    RECT 22.7 88.02 22.98 88.78 ;
    RECT 22.7 87.26 22.98 88.02 ;
    RECT 22.7 86.5 22.98 87.26 ;
    RECT 22.7 85.74 22.98 86.5 ;
    RECT 22.7 84.98 22.98 85.74 ;
    RECT 22.7 84.22 22.98 84.98 ;
    RECT 22.7 83.46 22.98 84.22 ;
    RECT 22.7 82.7 22.98 83.46 ;
    RECT 22.7 81.94 22.98 82.7 ;
    RECT 22.7 81.18 22.98 81.94 ;
    RECT 22.7 80.42 22.98 81.18 ;
    RECT 22.7 79.66 22.98 80.42 ;
    RECT 22.7 78.9 22.98 79.66 ;
    RECT 22.7 78.14 22.98 78.9 ;
    RECT 22.7 77.38 22.98 78.14 ;
    RECT 22.7 76.62 22.98 77.38 ;
    RECT 22.7 75.86 22.98 76.62 ;
    RECT 22.7 75.1 22.98 75.86 ;
    RECT 22.7 74.34 22.98 75.1 ;
    RECT 22.7 73.58 22.98 74.34 ;
    RECT 22.7 72.82 22.98 73.58 ;
    RECT 22.7 72.06 22.98 72.82 ;
    RECT 22.7 71.3 22.98 72.06 ;
    RECT 22.7 70.54 22.98 71.3 ;
    RECT 22.7 69.78 22.98 70.54 ;
    RECT 22.7 69.02 22.98 69.78 ;
    RECT 22.7 68.26 22.98 69.02 ;
    RECT 22.7 67.5 22.98 68.26 ;
    RECT 22.7 66.74 22.98 67.5 ;
    RECT 22.7 65.98 22.98 66.74 ;
    RECT 22.7 65.22 22.98 65.98 ;
    RECT 22.7 64.46 22.98 65.22 ;
    RECT 22.7 63.7 22.98 64.46 ;
    RECT 22.7 62.94 22.98 63.7 ;
    RECT 22.7 108.54 22.98 109.3 ;
    RECT 22.7 62.18 22.98 62.94 ;
    RECT 22.7 61.42 22.98 62.18 ;
    RECT 22.7 60.66 22.98 61.42 ;
    RECT 22.7 59.92 22.98 60.66 ;
    RECT 22.7 59.16 22.98 59.92 ;
    RECT 22.7 58.4 22.98 59.16 ;
    RECT 22.7 57.64 22.98 58.4 ;
    RECT 22.7 56.88 22.98 57.64 ;
    RECT 22.7 56.12 22.98 56.88 ;
    RECT 22.7 55.36 22.98 56.12 ;
    RECT 22.7 16.6 22.98 17.36 ;
    RECT 22.7 15.84 22.98 16.6 ;
    RECT 22.7 15.08 22.98 15.84 ;
    RECT 22.7 14.32 22.98 15.08 ;
    RECT 22.7 13.56 22.98 14.32 ;
    RECT 22.7 12.8 22.98 13.56 ;
    RECT 22.7 12.04 22.98 12.8 ;
    RECT 22.7 9.81 22.98 11.28 ;
    RECT 22.7 54.6 22.98 55.36 ;
    RECT 22.7 53.84 22.98 54.6 ;
    RECT 22.7 53.08 22.98 53.84 ;
    RECT 22.7 52.32 22.98 53.08 ;
    RECT 22.7 51.56 22.98 52.32 ;
    RECT 22.7 50.8 22.98 51.56 ;
    RECT 22.7 50.04 22.98 50.8 ;
    RECT 22.7 49.28 22.98 50.04 ;
    RECT 22.7 48.52 22.98 49.28 ;
    RECT 22.7 47.76 22.98 48.52 ;
    RECT 22.7 11.28 22.98 12.04 ;
    RECT 22.7 47.0 22.98 47.76 ;
    RECT 22.7 46.24 22.98 47.0 ;
    RECT 22.7 45.48 22.98 46.24 ;
    RECT 22.7 44.72 22.98 45.48 ;
    RECT 22.7 43.96 22.98 44.72 ;
    RECT 22.7 43.2 22.98 43.96 ;
    RECT 22.7 42.44 22.98 43.2 ;
    RECT 22.7 41.68 22.98 42.44 ;
    RECT 22.7 40.92 22.98 41.68 ;
    RECT 22.7 40.16 22.98 40.92 ;
    RECT 22.7 109.3 22.98 110.77 ;
    RECT 22.7 39.4 22.98 40.16 ;
    RECT 22.7 38.64 22.98 39.4 ;
    RECT 22.7 37.88 22.98 38.64 ;
    RECT 22.7 37.12 22.98 37.88 ;
    RECT 22.7 36.36 22.98 37.12 ;
    RECT 22.7 35.6 22.98 36.36 ;
    RECT 22.7 34.84 22.98 35.6 ;
    RECT 22.7 34.08 22.98 34.84 ;
    RECT 22.7 107.78 22.98 108.54 ;
    RECT 22.7 33.32 22.98 34.08 ;
    RECT 22.7 107.02 22.98 107.78 ;
    RECT 22.7 32.56 22.98 33.32 ;
    RECT 22.7 106.26 22.98 107.02 ;
    RECT 22.7 105.5 22.98 106.26 ;
    RECT 22.7 104.74 22.98 105.5 ;
    RECT 22.7 103.98 22.98 104.74 ;
    RECT 22.7 103.22 22.98 103.98 ;
    RECT 22.7 102.46 22.98 103.22 ;
    RECT 22.7 101.7 22.98 102.46 ;
    RECT 22.7 100.94 22.98 101.7 ;
    RECT 1.0 31.8 1.28 32.56 ;
    RECT 1.0 31.04 1.28 31.8 ;
    RECT 1.0 30.28 1.28 31.04 ;
    RECT 1.0 29.52 1.28 30.28 ;
    RECT 1.0 28.76 1.28 29.52 ;
    RECT 1.0 28.0 1.28 28.76 ;
    RECT 1.0 27.24 1.28 28.0 ;
    RECT 1.0 26.48 1.28 27.24 ;
    RECT 1.0 100.18 1.28 100.94 ;
    RECT 1.0 25.72 1.28 26.48 ;
    RECT 1.0 99.42 1.28 100.18 ;
    RECT 1.0 24.96 1.28 25.72 ;
    RECT 1.0 98.66 1.28 99.42 ;
    RECT 1.0 97.9 1.28 98.66 ;
    RECT 1.0 97.14 1.28 97.9 ;
    RECT 1.0 96.38 1.28 97.14 ;
    RECT 1.0 95.62 1.28 96.38 ;
    RECT 1.0 94.86 1.28 95.62 ;
    RECT 1.0 94.1 1.28 94.86 ;
    RECT 1.0 93.34 1.28 94.1 ;
    RECT 1.0 24.2 1.28 24.96 ;
    RECT 1.0 23.44 1.28 24.2 ;
    RECT 1.0 22.68 1.28 23.44 ;
    RECT 1.0 21.92 1.28 22.68 ;
    RECT 1.0 21.16 1.28 21.92 ;
    RECT 1.0 20.4 1.28 21.16 ;
    RECT 1.0 19.64 1.28 20.4 ;
    RECT 1.0 18.88 1.28 19.64 ;
    RECT 1.0 92.58 1.28 93.34 ;
    RECT 1.0 18.12 1.28 18.88 ;
    RECT 1.0 91.82 1.28 92.58 ;
    RECT 1.0 17.36 1.28 18.12 ;
    RECT 1.0 91.06 1.28 91.82 ;
    RECT 1.0 90.3 1.28 91.06 ;
    RECT 1.0 89.54 1.28 90.3 ;
    RECT 1.0 88.78 1.28 89.54 ;
    RECT 1.0 88.02 1.28 88.78 ;
    RECT 1.0 87.26 1.28 88.02 ;
    RECT 1.0 86.5 1.28 87.26 ;
    RECT 1.0 85.74 1.28 86.5 ;
    RECT 1.0 84.98 1.28 85.74 ;
    RECT 1.0 84.22 1.28 84.98 ;
    RECT 1.0 83.46 1.28 84.22 ;
    RECT 1.0 82.7 1.28 83.46 ;
    RECT 1.0 81.94 1.28 82.7 ;
    RECT 1.0 81.18 1.28 81.94 ;
    RECT 1.0 80.42 1.28 81.18 ;
    RECT 1.0 79.66 1.28 80.42 ;
    RECT 1.0 78.9 1.28 79.66 ;
    RECT 1.0 78.14 1.28 78.9 ;
    RECT 1.0 77.38 1.28 78.14 ;
    RECT 1.0 76.62 1.28 77.38 ;
    RECT 1.0 75.86 1.28 76.62 ;
    RECT 1.0 75.1 1.28 75.86 ;
    RECT 1.0 74.34 1.28 75.1 ;
    RECT 1.0 73.58 1.28 74.34 ;
    RECT 1.0 72.82 1.28 73.58 ;
    RECT 1.0 72.06 1.28 72.82 ;
    RECT 1.0 71.3 1.28 72.06 ;
    RECT 1.0 70.54 1.28 71.3 ;
    RECT 1.0 69.78 1.28 70.54 ;
    RECT 1.0 69.02 1.28 69.78 ;
    RECT 1.0 68.26 1.28 69.02 ;
    RECT 1.0 67.5 1.28 68.26 ;
    RECT 1.0 66.74 1.28 67.5 ;
    RECT 1.0 65.98 1.28 66.74 ;
    RECT 1.0 65.22 1.28 65.98 ;
    RECT 1.0 64.46 1.28 65.22 ;
    RECT 1.0 63.7 1.28 64.46 ;
    RECT 1.0 62.94 1.28 63.7 ;
    RECT 1.0 108.54 1.28 109.3 ;
    RECT 1.0 62.18 1.28 62.94 ;
    RECT 1.0 61.42 1.28 62.18 ;
    RECT 1.0 60.66 1.28 61.42 ;
    RECT 1.0 59.92 1.28 60.66 ;
    RECT 1.0 59.16 1.28 59.92 ;
    RECT 1.0 58.4 1.28 59.16 ;
    RECT 1.0 57.64 1.28 58.4 ;
    RECT 1.0 56.88 1.28 57.64 ;
    RECT 1.0 56.12 1.28 56.88 ;
    RECT 1.0 55.36 1.28 56.12 ;
    RECT 1.0 16.6 1.28 17.36 ;
    RECT 1.0 15.84 1.28 16.6 ;
    RECT 1.0 15.08 1.28 15.84 ;
    RECT 1.0 14.32 1.28 15.08 ;
    RECT 1.0 13.56 1.28 14.32 ;
    RECT 1.0 12.8 1.28 13.56 ;
    RECT 1.0 12.04 1.28 12.8 ;
    RECT 1.0 9.81 1.28 11.28 ;
    RECT 1.0 54.6 1.28 55.36 ;
    RECT 1.0 53.84 1.28 54.6 ;
    RECT 1.0 53.08 1.28 53.84 ;
    RECT 1.0 52.32 1.28 53.08 ;
    RECT 1.0 51.56 1.28 52.32 ;
    RECT 1.0 50.8 1.28 51.56 ;
    RECT 1.0 50.04 1.28 50.8 ;
    RECT 1.0 49.28 1.28 50.04 ;
    RECT 1.0 48.52 1.28 49.28 ;
    RECT 1.0 47.76 1.28 48.52 ;
    RECT 1.0 11.28 1.28 12.04 ;
    RECT 1.0 47.0 1.28 47.76 ;
    RECT 1.0 46.24 1.28 47.0 ;
    RECT 1.0 45.48 1.28 46.24 ;
    RECT 1.0 44.72 1.28 45.48 ;
    RECT 1.0 43.96 1.28 44.72 ;
    RECT 1.0 43.2 1.28 43.96 ;
    RECT 1.0 42.44 1.28 43.2 ;
    RECT 1.0 41.68 1.28 42.44 ;
    RECT 1.0 40.92 1.28 41.68 ;
    RECT 1.0 40.16 1.28 40.92 ;
    RECT 1.0 109.3 1.28 110.77 ;
    RECT 1.0 39.4 1.28 40.16 ;
    RECT 1.0 38.64 1.28 39.4 ;
    RECT 1.0 37.88 1.28 38.64 ;
    RECT 1.0 37.12 1.28 37.88 ;
    RECT 1.0 36.36 1.28 37.12 ;
    RECT 1.0 35.6 1.28 36.36 ;
    RECT 1.0 34.84 1.28 35.6 ;
    RECT 1.0 34.08 1.28 34.84 ;
    RECT 1.0 107.78 1.28 108.54 ;
    RECT 1.0 33.32 1.28 34.08 ;
    RECT 1.0 107.02 1.28 107.78 ;
    RECT 1.0 32.56 1.28 33.32 ;
    RECT 1.0 106.26 1.28 107.02 ;
    RECT 1.0 105.5 1.28 106.26 ;
    RECT 1.0 104.74 1.28 105.5 ;
    RECT 1.0 103.98 1.28 104.74 ;
    RECT 1.0 103.22 1.28 103.98 ;
    RECT 1.0 102.46 1.28 103.22 ;
    RECT 1.0 101.7 1.28 102.46 ;
    RECT 1.0 100.94 1.28 101.7 ;
    RECT 16.5 0.43 16.78 0.78 ;
    RECT 13.4 0.43 13.68 0.78 ;
    RECT 22.7 0.43 22.98 0.78 ;
    RECT 19.6 0.43 19.88 0.78 ;
    RECT 4.1 0.43 4.38 0.78 ;
    RECT 1.0 0.43 1.28 0.78 ;
    RECT 10.3 0.43 10.58 0.78 ;
    RECT 7.2 0.43 7.48 0.78 ;
    RECT 22.7 1.32 22.98 2.76 ;
    RECT 19.6 1.32 19.88 2.76 ;
    RECT 10.3 1.32 10.58 2.76 ;
    RECT 7.2 1.32 7.48 2.76 ;
    RECT 16.5 1.32 16.78 2.76 ;
    RECT 13.4 1.32 13.68 2.76 ;
    RECT 4.1 1.32 4.38 2.76 ;
    RECT 1.0 1.32 1.28 2.76 ;
    RECT 22.7 2.76 22.98 9.81 ;
    RECT 19.6 2.76 19.88 9.81 ;
    RECT 4.1 2.76 4.38 9.81 ;
    RECT 1.0 2.76 1.28 9.81 ;
    RECT 10.3 2.76 10.58 9.81 ;
    RECT 7.2 2.76 7.48 9.81 ;
    RECT 16.5 2.76 16.78 9.81 ;
    RECT 13.4 2.76 13.68 9.81 ;
    RECT 10.3 0.78 10.58 1.32 ;
    RECT 7.2 0.78 7.48 1.32 ;
    RECT 16.5 0.78 16.78 1.32 ;
    RECT 13.4 0.78 13.68 1.32 ;
    RECT 22.7 0.78 22.98 1.32 ;
    RECT 19.6 0.78 19.88 1.32 ;
    RECT 4.1 0.78 4.38 1.32 ;
    RECT 1.0 0.78 1.28 1.32 ;
    RECT 93.435 0.43 93.715 0.78 ;
    RECT 96.535 0.43 96.815 0.78 ;
    RECT 87.235 0.43 87.515 0.78 ;
    RECT 90.335 0.43 90.615 0.78 ;
    RECT 105.835 0.43 106.115 0.78 ;
    RECT 108.935 0.43 109.215 0.78 ;
    RECT 99.635 0.43 99.915 0.78 ;
    RECT 102.735 0.43 103.015 0.78 ;
    RECT 87.235 1.32 87.515 2.76 ;
    RECT 90.335 1.32 90.615 2.76 ;
    RECT 99.635 1.32 99.915 2.76 ;
    RECT 102.735 1.32 103.015 2.76 ;
    RECT 93.435 1.32 93.715 2.76 ;
    RECT 96.535 1.32 96.815 2.76 ;
    RECT 105.835 1.32 106.115 2.76 ;
    RECT 108.935 1.32 109.215 2.76 ;
    RECT 87.235 2.76 87.515 9.81 ;
    RECT 90.335 2.76 90.615 9.81 ;
    RECT 105.835 2.76 106.115 9.81 ;
    RECT 108.935 2.76 109.215 9.81 ;
    RECT 99.635 2.76 99.915 9.81 ;
    RECT 102.735 2.76 103.015 9.81 ;
    RECT 93.435 2.76 93.715 9.81 ;
    RECT 96.535 2.76 96.815 9.81 ;
    RECT 99.635 0.78 99.915 1.32 ;
    RECT 102.735 0.78 103.015 1.32 ;
    RECT 93.435 0.78 93.715 1.32 ;
    RECT 96.535 0.78 96.815 1.32 ;
    RECT 87.235 0.78 87.515 1.32 ;
    RECT 90.335 0.78 90.615 1.32 ;
    RECT 105.835 0.78 106.115 1.32 ;
    RECT 108.935 0.78 109.215 1.32 ;
    #obstructions of filtered out pwrgnd shapes
    RECT 76.07 0.43 76.17 0.78 ;
    RECT 76.765 0.43 76.865 0.78 ;
    RECT 53.69 1.865 53.83 9.485 ;
    RECT 74.67 0.78 74.77 1.235 ;
    RECT 76.07 110.77 76.17 111.055 ;
    RECT 76.765 110.77 76.865 111.055 ;
    END
  END rf_2p_hde

END LIBRARY

